/* ******************************** */
/* Arithmetic Module Generator	*/
/* Carry Propagate Array Multiplier */
/* Multiplier Size: 16 */
/* Inputs: a[15 :0], b[15 :0] */
/* Output: m[31 :0] */
/* ******************************** */

`timescale 1ns/10ps 

module HA (I1, I2, sum, carry);
input I1, I2;
output sum, carry;
xor (sum, I1, I2);
and (carry, I1, I2);
endmodule

module FA (I1, I2, I3, sum, carry);
input I1, I2, I3;
output sum, carry;

wire xout,o1,o2;
xor (xout, I1, I2);
xor (sum, xout, I3);
and (o1, I1, I2);
and (o2, xout, I3);
or (carry, o1, o2);
endmodule

module multiplier (a, b, m);
input	[15 :0] a;
input	[15 :0] b;
output	[31 :0] m;

wire	[255 :1]	pp;
wire	[14 :0]	r1c;
wire	[14 :1]	r1s;
wire	[14 :0]	r2c;
wire	[14 :1]	r2s;
wire	[14 :0]	r3c;
wire	[14 :1]	r3s;
wire	[14 :0]	r4c;
wire	[14 :1]	r4s;
wire	[14 :0]	r5c;
wire	[14 :1]	r5s;
wire	[14 :0]	r6c;
wire	[14 :1]	r6s;
wire	[14 :0]	r7c;
wire	[14 :1]	r7s;
wire	[14 :0]	r8c;
wire	[14 :1]	r8s;
wire	[14 :0]	r9c;
wire	[14 :1]	r9s;
wire	[14 :0]	r10c;
wire	[14 :1]	r10s;
wire	[14 :0]	r11c;
wire	[14 :1]	r11s;
wire	[14 :0]	r12c;
wire	[14 :1]	r12s;
wire	[14 :0]	r13c;
wire	[14 :1]	r13s;
wire	[14 :0]	r14c;
wire	[14 :1]	r14s;
wire	[14 :0]	r15c;
wire	[14 :1]	r15s;
wire	[13 :0]	r16c;

and	(m[0], a[0], b[0]);
and	(pp[1], a[0], b[1]);
and	(pp[2], a[0], b[2]);
and	(pp[3], a[0], b[3]);
and	(pp[4], a[0], b[4]);
and	(pp[5], a[0], b[5]);
and	(pp[6], a[0], b[6]);
and	(pp[7], a[0], b[7]);
and	(pp[8], a[0], b[8]);
and	(pp[9], a[0], b[9]);
and	(pp[10], a[0], b[10]);
and	(pp[11], a[0], b[11]);
and	(pp[12], a[0], b[12]);
and	(pp[13], a[0], b[13]);
and	(pp[14], a[0], b[14]);
and	(pp[15], a[0], b[15]);
and	(pp[16], a[1], b[0]);
and	(pp[17], a[1], b[1]);
and	(pp[18], a[1], b[2]);
and	(pp[19], a[1], b[3]);
and	(pp[20], a[1], b[4]);
and	(pp[21], a[1], b[5]);
and	(pp[22], a[1], b[6]);
and	(pp[23], a[1], b[7]);
and	(pp[24], a[1], b[8]);
and	(pp[25], a[1], b[9]);
and	(pp[26], a[1], b[10]);
and	(pp[27], a[1], b[11]);
and	(pp[28], a[1], b[12]);
and	(pp[29], a[1], b[13]);
and	(pp[30], a[1], b[14]);
and	(pp[31], a[1], b[15]);
and	(pp[32], a[2], b[0]);
and	(pp[33], a[2], b[1]);
and	(pp[34], a[2], b[2]);
and	(pp[35], a[2], b[3]);
and	(pp[36], a[2], b[4]);
and	(pp[37], a[2], b[5]);
and	(pp[38], a[2], b[6]);
and	(pp[39], a[2], b[7]);
and	(pp[40], a[2], b[8]);
and	(pp[41], a[2], b[9]);
and	(pp[42], a[2], b[10]);
and	(pp[43], a[2], b[11]);
and	(pp[44], a[2], b[12]);
and	(pp[45], a[2], b[13]);
and	(pp[46], a[2], b[14]);
and	(pp[47], a[2], b[15]);
and	(pp[48], a[3], b[0]);
and	(pp[49], a[3], b[1]);
and	(pp[50], a[3], b[2]);
and	(pp[51], a[3], b[3]);
and	(pp[52], a[3], b[4]);
and	(pp[53], a[3], b[5]);
and	(pp[54], a[3], b[6]);
and	(pp[55], a[3], b[7]);
and	(pp[56], a[3], b[8]);
and	(pp[57], a[3], b[9]);
and	(pp[58], a[3], b[10]);
and	(pp[59], a[3], b[11]);
and	(pp[60], a[3], b[12]);
and	(pp[61], a[3], b[13]);
and	(pp[62], a[3], b[14]);
and	(pp[63], a[3], b[15]);
and	(pp[64], a[4], b[0]);
and	(pp[65], a[4], b[1]);
and	(pp[66], a[4], b[2]);
and	(pp[67], a[4], b[3]);
and	(pp[68], a[4], b[4]);
and	(pp[69], a[4], b[5]);
and	(pp[70], a[4], b[6]);
and	(pp[71], a[4], b[7]);
and	(pp[72], a[4], b[8]);
and	(pp[73], a[4], b[9]);
and	(pp[74], a[4], b[10]);
and	(pp[75], a[4], b[11]);
and	(pp[76], a[4], b[12]);
and	(pp[77], a[4], b[13]);
and	(pp[78], a[4], b[14]);
and	(pp[79], a[4], b[15]);
and	(pp[80], a[5], b[0]);
and	(pp[81], a[5], b[1]);
and	(pp[82], a[5], b[2]);
and	(pp[83], a[5], b[3]);
and	(pp[84], a[5], b[4]);
and	(pp[85], a[5], b[5]);
and	(pp[86], a[5], b[6]);
and	(pp[87], a[5], b[7]);
and	(pp[88], a[5], b[8]);
and	(pp[89], a[5], b[9]);
and	(pp[90], a[5], b[10]);
and	(pp[91], a[5], b[11]);
and	(pp[92], a[5], b[12]);
and	(pp[93], a[5], b[13]);
and	(pp[94], a[5], b[14]);
and	(pp[95], a[5], b[15]);
and	(pp[96], a[6], b[0]);
and	(pp[97], a[6], b[1]);
and	(pp[98], a[6], b[2]);
and	(pp[99], a[6], b[3]);
and	(pp[100], a[6], b[4]);
and	(pp[101], a[6], b[5]);
and	(pp[102], a[6], b[6]);
and	(pp[103], a[6], b[7]);
and	(pp[104], a[6], b[8]);
and	(pp[105], a[6], b[9]);
and	(pp[106], a[6], b[10]);
and	(pp[107], a[6], b[11]);
and	(pp[108], a[6], b[12]);
and	(pp[109], a[6], b[13]);
and	(pp[110], a[6], b[14]);
and	(pp[111], a[6], b[15]);
and	(pp[112], a[7], b[0]);
and	(pp[113], a[7], b[1]);
and	(pp[114], a[7], b[2]);
and	(pp[115], a[7], b[3]);
and	(pp[116], a[7], b[4]);
and	(pp[117], a[7], b[5]);
and	(pp[118], a[7], b[6]);
and	(pp[119], a[7], b[7]);
and	(pp[120], a[7], b[8]);
and	(pp[121], a[7], b[9]);
and	(pp[122], a[7], b[10]);
and	(pp[123], a[7], b[11]);
and	(pp[124], a[7], b[12]);
and	(pp[125], a[7], b[13]);
and	(pp[126], a[7], b[14]);
and	(pp[127], a[7], b[15]);
and	(pp[128], a[8], b[0]);
and	(pp[129], a[8], b[1]);
and	(pp[130], a[8], b[2]);
and	(pp[131], a[8], b[3]);
and	(pp[132], a[8], b[4]);
and	(pp[133], a[8], b[5]);
and	(pp[134], a[8], b[6]);
and	(pp[135], a[8], b[7]);
and	(pp[136], a[8], b[8]);
and	(pp[137], a[8], b[9]);
and	(pp[138], a[8], b[10]);
and	(pp[139], a[8], b[11]);
and	(pp[140], a[8], b[12]);
and	(pp[141], a[8], b[13]);
and	(pp[142], a[8], b[14]);
and	(pp[143], a[8], b[15]);
and	(pp[144], a[9], b[0]);
and	(pp[145], a[9], b[1]);
and	(pp[146], a[9], b[2]);
and	(pp[147], a[9], b[3]);
and	(pp[148], a[9], b[4]);
and	(pp[149], a[9], b[5]);
and	(pp[150], a[9], b[6]);
and	(pp[151], a[9], b[7]);
and	(pp[152], a[9], b[8]);
and	(pp[153], a[9], b[9]);
and	(pp[154], a[9], b[10]);
and	(pp[155], a[9], b[11]);
and	(pp[156], a[9], b[12]);
and	(pp[157], a[9], b[13]);
and	(pp[158], a[9], b[14]);
and	(pp[159], a[9], b[15]);
and	(pp[160], a[10], b[0]);
and	(pp[161], a[10], b[1]);
and	(pp[162], a[10], b[2]);
and	(pp[163], a[10], b[3]);
and	(pp[164], a[10], b[4]);
and	(pp[165], a[10], b[5]);
and	(pp[166], a[10], b[6]);
and	(pp[167], a[10], b[7]);
and	(pp[168], a[10], b[8]);
and	(pp[169], a[10], b[9]);
and	(pp[170], a[10], b[10]);
and	(pp[171], a[10], b[11]);
and	(pp[172], a[10], b[12]);
and	(pp[173], a[10], b[13]);
and	(pp[174], a[10], b[14]);
and	(pp[175], a[10], b[15]);
and	(pp[176], a[11], b[0]);
and	(pp[177], a[11], b[1]);
and	(pp[178], a[11], b[2]);
and	(pp[179], a[11], b[3]);
and	(pp[180], a[11], b[4]);
and	(pp[181], a[11], b[5]);
and	(pp[182], a[11], b[6]);
and	(pp[183], a[11], b[7]);
and	(pp[184], a[11], b[8]);
and	(pp[185], a[11], b[9]);
and	(pp[186], a[11], b[10]);
and	(pp[187], a[11], b[11]);
and	(pp[188], a[11], b[12]);
and	(pp[189], a[11], b[13]);
and	(pp[190], a[11], b[14]);
and	(pp[191], a[11], b[15]);
and	(pp[192], a[12], b[0]);
and	(pp[193], a[12], b[1]);
and	(pp[194], a[12], b[2]);
and	(pp[195], a[12], b[3]);
and	(pp[196], a[12], b[4]);
and	(pp[197], a[12], b[5]);
and	(pp[198], a[12], b[6]);
and	(pp[199], a[12], b[7]);
and	(pp[200], a[12], b[8]);
and	(pp[201], a[12], b[9]);
and	(pp[202], a[12], b[10]);
and	(pp[203], a[12], b[11]);
and	(pp[204], a[12], b[12]);
and	(pp[205], a[12], b[13]);
and	(pp[206], a[12], b[14]);
and	(pp[207], a[12], b[15]);
and	(pp[208], a[13], b[0]);
and	(pp[209], a[13], b[1]);
and	(pp[210], a[13], b[2]);
and	(pp[211], a[13], b[3]);
and	(pp[212], a[13], b[4]);
and	(pp[213], a[13], b[5]);
and	(pp[214], a[13], b[6]);
and	(pp[215], a[13], b[7]);
and	(pp[216], a[13], b[8]);
and	(pp[217], a[13], b[9]);
and	(pp[218], a[13], b[10]);
and	(pp[219], a[13], b[11]);
and	(pp[220], a[13], b[12]);
and	(pp[221], a[13], b[13]);
and	(pp[222], a[13], b[14]);
and	(pp[223], a[13], b[15]);
and	(pp[224], a[14], b[0]);
and	(pp[225], a[14], b[1]);
and	(pp[226], a[14], b[2]);
and	(pp[227], a[14], b[3]);
and	(pp[228], a[14], b[4]);
and	(pp[229], a[14], b[5]);
and	(pp[230], a[14], b[6]);
and	(pp[231], a[14], b[7]);
and	(pp[232], a[14], b[8]);
and	(pp[233], a[14], b[9]);
and	(pp[234], a[14], b[10]);
and	(pp[235], a[14], b[11]);
and	(pp[236], a[14], b[12]);
and	(pp[237], a[14], b[13]);
and	(pp[238], a[14], b[14]);
and	(pp[239], a[14], b[15]);
and	(pp[240], a[15], b[0]);
and	(pp[241], a[15], b[1]);
and	(pp[242], a[15], b[2]);
and	(pp[243], a[15], b[3]);
and	(pp[244], a[15], b[4]);
and	(pp[245], a[15], b[5]);
and	(pp[246], a[15], b[6]);
and	(pp[247], a[15], b[7]);
and	(pp[248], a[15], b[8]);
and	(pp[249], a[15], b[9]);
and	(pp[250], a[15], b[10]);
and	(pp[251], a[15], b[11]);
and	(pp[252], a[15], b[12]);
and	(pp[253], a[15], b[13]);
and	(pp[254], a[15], b[14]);
and	(pp[255], a[15], b[15]);

HA	inst257	(pp[16], pp[1], m[1], r1c[0]);
FA	inst258	(pp[17], pp[2], r1c[0], r1s[1], r1c[1]);
FA	inst259	(pp[18], pp[3], r1c[1], r1s[2], r1c[2]);
FA	inst260	(pp[19], pp[4], r1c[2], r1s[3], r1c[3]);
FA	inst261	(pp[20], pp[5], r1c[3], r1s[4], r1c[4]);
FA	inst262	(pp[21], pp[6], r1c[4], r1s[5], r1c[5]);
FA	inst263	(pp[22], pp[7], r1c[5], r1s[6], r1c[6]);
FA	inst264	(pp[23], pp[8], r1c[6], r1s[7], r1c[7]);
FA	inst265	(pp[24], pp[9], r1c[7], r1s[8], r1c[8]);
FA	inst266	(pp[25], pp[10], r1c[8], r1s[9], r1c[9]);
FA	inst267	(pp[26], pp[11], r1c[9], r1s[10], r1c[10]);
FA	inst268	(pp[27], pp[12], r1c[10], r1s[11], r1c[11]);
FA	inst269	(pp[28], pp[13], r1c[11], r1s[12], r1c[12]);
FA	inst270	(pp[29], pp[14], r1c[12], r1s[13], r1c[13]);
FA	inst271	(pp[30], pp[15], r1c[13], r1s[14], r1c[14]);

HA	inst272	(r1s[1], pp[32], m[2], r2c[0]);
FA	inst273	(r1s[2], pp[33], r2c[0], r2s[1], r2c[1]);
FA	inst274	(r1s[3], pp[34], r2c[1], r2s[2], r2c[2]);
FA	inst275	(r1s[4], pp[35], r2c[2], r2s[3], r2c[3]);
FA	inst276	(r1s[5], pp[36], r2c[3], r2s[4], r2c[4]);
FA	inst277	(r1s[6], pp[37], r2c[4], r2s[5], r2c[5]);
FA	inst278	(r1s[7], pp[38], r2c[5], r2s[6], r2c[6]);
FA	inst279	(r1s[8], pp[39], r2c[6], r2s[7], r2c[7]);
FA	inst280	(r1s[9], pp[40], r2c[7], r2s[8], r2c[8]);
FA	inst281	(r1s[10], pp[41], r2c[8], r2s[9], r2c[9]);
FA	inst282	(r1s[11], pp[42], r2c[9], r2s[10], r2c[10]);
FA	inst283	(r1s[12], pp[43], r2c[10], r2s[11], r2c[11]);
FA	inst284	(r1s[13], pp[44], r2c[11], r2s[12], r2c[12]);
FA	inst285	(r1s[14], pp[45], r2c[12], r2s[13], r2c[13]);
FA	inst286	(r1c[14], pp[31], r2c[13], r2s[14], r2c[14]);

HA	inst287	(r2s[1], pp[48], m[3], r3c[0]);
FA	inst288	(r2s[2], pp[49], r3c[0], r3s[1], r3c[1]);
FA	inst289	(r2s[3], pp[50], r3c[1], r3s[2], r3c[2]);
FA	inst290	(r2s[4], pp[51], r3c[2], r3s[3], r3c[3]);
FA	inst291	(r2s[5], pp[52], r3c[3], r3s[4], r3c[4]);
FA	inst292	(r2s[6], pp[53], r3c[4], r3s[5], r3c[5]);
FA	inst293	(r2s[7], pp[54], r3c[5], r3s[6], r3c[6]);
FA	inst294	(r2s[8], pp[55], r3c[6], r3s[7], r3c[7]);
FA	inst295	(r2s[9], pp[56], r3c[7], r3s[8], r3c[8]);
FA	inst296	(r2s[10], pp[57], r3c[8], r3s[9], r3c[9]);
FA	inst297	(r2s[11], pp[58], r3c[9], r3s[10], r3c[10]);
FA	inst298	(r2s[12], pp[59], r3c[10], r3s[11], r3c[11]);
FA	inst299	(r2s[13], pp[60], r3c[11], r3s[12], r3c[12]);
FA	inst300	(r2s[14], pp[46], r3c[12], r3s[13], r3c[13]);
FA	inst301	(r2c[14], pp[47], r3c[13], r3s[14], r3c[14]);

HA	inst302	(r3s[1], pp[64], m[4], r4c[0]);
FA	inst303	(r3s[2], pp[65], r4c[0], r4s[1], r4c[1]);
FA	inst304	(r3s[3], pp[66], r4c[1], r4s[2], r4c[2]);
FA	inst305	(r3s[4], pp[67], r4c[2], r4s[3], r4c[3]);
FA	inst306	(r3s[5], pp[68], r4c[3], r4s[4], r4c[4]);
FA	inst307	(r3s[6], pp[69], r4c[4], r4s[5], r4c[5]);
FA	inst308	(r3s[7], pp[70], r4c[5], r4s[6], r4c[6]);
FA	inst309	(r3s[8], pp[71], r4c[6], r4s[7], r4c[7]);
FA	inst310	(r3s[9], pp[72], r4c[7], r4s[8], r4c[8]);
FA	inst311	(r3s[10], pp[73], r4c[8], r4s[9], r4c[9]);
FA	inst312	(r3s[11], pp[74], r4c[9], r4s[10], r4c[10]);
FA	inst313	(r3s[12], pp[75], r4c[10], r4s[11], r4c[11]);
FA	inst314	(r3s[13], pp[61], r4c[11], r4s[12], r4c[12]);
FA	inst315	(r3s[14], pp[62], r4c[12], r4s[13], r4c[13]);
FA	inst316	(r3c[14], pp[63], r4c[13], r4s[14], r4c[14]);

HA	inst317	(r4s[1], pp[80], m[5], r5c[0]);
FA	inst318	(r4s[2], pp[81], r5c[0], r5s[1], r5c[1]);
FA	inst319	(r4s[3], pp[82], r5c[1], r5s[2], r5c[2]);
FA	inst320	(r4s[4], pp[83], r5c[2], r5s[3], r5c[3]);
FA	inst321	(r4s[5], pp[84], r5c[3], r5s[4], r5c[4]);
FA	inst322	(r4s[6], pp[85], r5c[4], r5s[5], r5c[5]);
FA	inst323	(r4s[7], pp[86], r5c[5], r5s[6], r5c[6]);
FA	inst324	(r4s[8], pp[87], r5c[6], r5s[7], r5c[7]);
FA	inst325	(r4s[9], pp[88], r5c[7], r5s[8], r5c[8]);
FA	inst326	(r4s[10], pp[89], r5c[8], r5s[9], r5c[9]);
FA	inst327	(r4s[11], pp[90], r5c[9], r5s[10], r5c[10]);
FA	inst328	(r4s[12], pp[76], r5c[10], r5s[11], r5c[11]);
FA	inst329	(r4s[13], pp[77], r5c[11], r5s[12], r5c[12]);
FA	inst330	(r4s[14], pp[78], r5c[12], r5s[13], r5c[13]);
FA	inst331	(r4c[14], pp[79], r5c[13], r5s[14], r5c[14]);

HA	inst332	(r5s[1], pp[96], m[6], r6c[0]);
FA	inst333	(r5s[2], pp[97], r6c[0], r6s[1], r6c[1]);
FA	inst334	(r5s[3], pp[98], r6c[1], r6s[2], r6c[2]);
FA	inst335	(r5s[4], pp[99], r6c[2], r6s[3], r6c[3]);
FA	inst336	(r5s[5], pp[100], r6c[3], r6s[4], r6c[4]);
FA	inst337	(r5s[6], pp[101], r6c[4], r6s[5], r6c[5]);
FA	inst338	(r5s[7], pp[102], r6c[5], r6s[6], r6c[6]);
FA	inst339	(r5s[8], pp[103], r6c[6], r6s[7], r6c[7]);
FA	inst340	(r5s[9], pp[104], r6c[7], r6s[8], r6c[8]);
FA	inst341	(r5s[10], pp[105], r6c[8], r6s[9], r6c[9]);
FA	inst342	(r5s[11], pp[91], r6c[9], r6s[10], r6c[10]);
FA	inst343	(r5s[12], pp[92], r6c[10], r6s[11], r6c[11]);
FA	inst344	(r5s[13], pp[93], r6c[11], r6s[12], r6c[12]);
FA	inst345	(r5s[14], pp[94], r6c[12], r6s[13], r6c[13]);
FA	inst346	(r5c[14], pp[95], r6c[13], r6s[14], r6c[14]);

HA	inst347	(r6s[1], pp[112], m[7], r7c[0]);
FA	inst348	(r6s[2], pp[113], r7c[0], r7s[1], r7c[1]);
FA	inst349	(r6s[3], pp[114], r7c[1], r7s[2], r7c[2]);
FA	inst350	(r6s[4], pp[115], r7c[2], r7s[3], r7c[3]);
FA	inst351	(r6s[5], pp[116], r7c[3], r7s[4], r7c[4]);
FA	inst352	(r6s[6], pp[117], r7c[4], r7s[5], r7c[5]);
FA	inst353	(r6s[7], pp[118], r7c[5], r7s[6], r7c[6]);
FA	inst354	(r6s[8], pp[119], r7c[6], r7s[7], r7c[7]);
FA	inst355	(r6s[9], pp[120], r7c[7], r7s[8], r7c[8]);
FA	inst356	(r6s[10], pp[106], r7c[8], r7s[9], r7c[9]);
FA	inst357	(r6s[11], pp[107], r7c[9], r7s[10], r7c[10]);
FA	inst358	(r6s[12], pp[108], r7c[10], r7s[11], r7c[11]);
FA	inst359	(r6s[13], pp[109], r7c[11], r7s[12], r7c[12]);
FA	inst360	(r6s[14], pp[110], r7c[12], r7s[13], r7c[13]);
FA	inst361	(r6c[14], pp[111], r7c[13], r7s[14], r7c[14]);

HA	inst362	(r7s[1], pp[128], m[8], r8c[0]);
FA	inst363	(r7s[2], pp[129], r8c[0], r8s[1], r8c[1]);
FA	inst364	(r7s[3], pp[130], r8c[1], r8s[2], r8c[2]);
FA	inst365	(r7s[4], pp[131], r8c[2], r8s[3], r8c[3]);
FA	inst366	(r7s[5], pp[132], r8c[3], r8s[4], r8c[4]);
FA	inst367	(r7s[6], pp[133], r8c[4], r8s[5], r8c[5]);
FA	inst368	(r7s[7], pp[134], r8c[5], r8s[6], r8c[6]);
FA	inst369	(r7s[8], pp[135], r8c[6], r8s[7], r8c[7]);
FA	inst370	(r7s[9], pp[121], r8c[7], r8s[8], r8c[8]);
FA	inst371	(r7s[10], pp[122], r8c[8], r8s[9], r8c[9]);
FA	inst372	(r7s[11], pp[123], r8c[9], r8s[10], r8c[10]);
FA	inst373	(r7s[12], pp[124], r8c[10], r8s[11], r8c[11]);
FA	inst374	(r7s[13], pp[125], r8c[11], r8s[12], r8c[12]);
FA	inst375	(r7s[14], pp[126], r8c[12], r8s[13], r8c[13]);
FA	inst376	(r7c[14], pp[127], r8c[13], r8s[14], r8c[14]);

HA	inst377	(r8s[1], pp[144], m[9], r9c[0]);
FA	inst378	(r8s[2], pp[145], r9c[0], r9s[1], r9c[1]);
FA	inst379	(r8s[3], pp[146], r9c[1], r9s[2], r9c[2]);
FA	inst380	(r8s[4], pp[147], r9c[2], r9s[3], r9c[3]);
FA	inst381	(r8s[5], pp[148], r9c[3], r9s[4], r9c[4]);
FA	inst382	(r8s[6], pp[149], r9c[4], r9s[5], r9c[5]);
FA	inst383	(r8s[7], pp[150], r9c[5], r9s[6], r9c[6]);
FA	inst384	(r8s[8], pp[136], r9c[6], r9s[7], r9c[7]);
FA	inst385	(r8s[9], pp[137], r9c[7], r9s[8], r9c[8]);
FA	inst386	(r8s[10], pp[138], r9c[8], r9s[9], r9c[9]);
FA	inst387	(r8s[11], pp[139], r9c[9], r9s[10], r9c[10]);
FA	inst388	(r8s[12], pp[140], r9c[10], r9s[11], r9c[11]);
FA	inst389	(r8s[13], pp[141], r9c[11], r9s[12], r9c[12]);
FA	inst390	(r8s[14], pp[142], r9c[12], r9s[13], r9c[13]);
FA	inst391	(r8c[14], pp[143], r9c[13], r9s[14], r9c[14]);

HA	inst392	(r9s[1], pp[160], m[10], r10c[0]);
FA	inst393	(r9s[2], pp[161], r10c[0], r10s[1], r10c[1]);
FA	inst394	(r9s[3], pp[162], r10c[1], r10s[2], r10c[2]);
FA	inst395	(r9s[4], pp[163], r10c[2], r10s[3], r10c[3]);
FA	inst396	(r9s[5], pp[164], r10c[3], r10s[4], r10c[4]);
FA	inst397	(r9s[6], pp[165], r10c[4], r10s[5], r10c[5]);
FA	inst398	(r9s[7], pp[151], r10c[5], r10s[6], r10c[6]);
FA	inst399	(r9s[8], pp[152], r10c[6], r10s[7], r10c[7]);
FA	inst400	(r9s[9], pp[153], r10c[7], r10s[8], r10c[8]);
FA	inst401	(r9s[10], pp[154], r10c[8], r10s[9], r10c[9]);
FA	inst402	(r9s[11], pp[155], r10c[9], r10s[10], r10c[10]);
FA	inst403	(r9s[12], pp[156], r10c[10], r10s[11], r10c[11]);
FA	inst404	(r9s[13], pp[157], r10c[11], r10s[12], r10c[12]);
FA	inst405	(r9s[14], pp[158], r10c[12], r10s[13], r10c[13]);
FA	inst406	(r9c[14], pp[159], r10c[13], r10s[14], r10c[14]);

HA	inst407	(r10s[1], pp[176], m[11], r11c[0]);
FA	inst408	(r10s[2], pp[177], r11c[0], r11s[1], r11c[1]);
FA	inst409	(r10s[3], pp[178], r11c[1], r11s[2], r11c[2]);
FA	inst410	(r10s[4], pp[179], r11c[2], r11s[3], r11c[3]);
FA	inst411	(r10s[5], pp[180], r11c[3], r11s[4], r11c[4]);
FA	inst412	(r10s[6], pp[166], r11c[4], r11s[5], r11c[5]);
FA	inst413	(r10s[7], pp[167], r11c[5], r11s[6], r11c[6]);
FA	inst414	(r10s[8], pp[168], r11c[6], r11s[7], r11c[7]);
FA	inst415	(r10s[9], pp[169], r11c[7], r11s[8], r11c[8]);
FA	inst416	(r10s[10], pp[170], r11c[8], r11s[9], r11c[9]);
FA	inst417	(r10s[11], pp[171], r11c[9], r11s[10], r11c[10]);
FA	inst418	(r10s[12], pp[172], r11c[10], r11s[11], r11c[11]);
FA	inst419	(r10s[13], pp[173], r11c[11], r11s[12], r11c[12]);
FA	inst420	(r10s[14], pp[174], r11c[12], r11s[13], r11c[13]);
FA	inst421	(r10c[14], pp[175], r11c[13], r11s[14], r11c[14]);

HA	inst422	(r11s[1], pp[192], m[12], r12c[0]);
FA	inst423	(r11s[2], pp[193], r12c[0], r12s[1], r12c[1]);
FA	inst424	(r11s[3], pp[194], r12c[1], r12s[2], r12c[2]);
FA	inst425	(r11s[4], pp[195], r12c[2], r12s[3], r12c[3]);
FA	inst426	(r11s[5], pp[181], r12c[3], r12s[4], r12c[4]);
FA	inst427	(r11s[6], pp[182], r12c[4], r12s[5], r12c[5]);
FA	inst428	(r11s[7], pp[183], r12c[5], r12s[6], r12c[6]);
FA	inst429	(r11s[8], pp[184], r12c[6], r12s[7], r12c[7]);
FA	inst430	(r11s[9], pp[185], r12c[7], r12s[8], r12c[8]);
FA	inst431	(r11s[10], pp[186], r12c[8], r12s[9], r12c[9]);
FA	inst432	(r11s[11], pp[187], r12c[9], r12s[10], r12c[10]);
FA	inst433	(r11s[12], pp[188], r12c[10], r12s[11], r12c[11]);
FA	inst434	(r11s[13], pp[189], r12c[11], r12s[12], r12c[12]);
FA	inst435	(r11s[14], pp[190], r12c[12], r12s[13], r12c[13]);
FA	inst436	(r11c[14], pp[191], r12c[13], r12s[14], r12c[14]);

HA	inst437	(r12s[1], pp[208], m[13], r13c[0]);
FA	inst438	(r12s[2], pp[209], r13c[0], r13s[1], r13c[1]);
FA	inst439	(r12s[3], pp[210], r13c[1], r13s[2], r13c[2]);
FA	inst440	(r12s[4], pp[196], r13c[2], r13s[3], r13c[3]);
FA	inst441	(r12s[5], pp[197], r13c[3], r13s[4], r13c[4]);
FA	inst442	(r12s[6], pp[198], r13c[4], r13s[5], r13c[5]);
FA	inst443	(r12s[7], pp[199], r13c[5], r13s[6], r13c[6]);
FA	inst444	(r12s[8], pp[200], r13c[6], r13s[7], r13c[7]);
FA	inst445	(r12s[9], pp[201], r13c[7], r13s[8], r13c[8]);
FA	inst446	(r12s[10], pp[202], r13c[8], r13s[9], r13c[9]);
FA	inst447	(r12s[11], pp[203], r13c[9], r13s[10], r13c[10]);
FA	inst448	(r12s[12], pp[204], r13c[10], r13s[11], r13c[11]);
FA	inst449	(r12s[13], pp[205], r13c[11], r13s[12], r13c[12]);
FA	inst450	(r12s[14], pp[206], r13c[12], r13s[13], r13c[13]);
FA	inst451	(r12c[14], pp[207], r13c[13], r13s[14], r13c[14]);

HA	inst452	(r13s[1], pp[224], m[14], r14c[0]);
FA	inst453	(r13s[2], pp[225], r14c[0], r14s[1], r14c[1]);
FA	inst454	(r13s[3], pp[211], r14c[1], r14s[2], r14c[2]);
FA	inst455	(r13s[4], pp[212], r14c[2], r14s[3], r14c[3]);
FA	inst456	(r13s[5], pp[213], r14c[3], r14s[4], r14c[4]);
FA	inst457	(r13s[6], pp[214], r14c[4], r14s[5], r14c[5]);
FA	inst458	(r13s[7], pp[215], r14c[5], r14s[6], r14c[6]);
FA	inst459	(r13s[8], pp[216], r14c[6], r14s[7], r14c[7]);
FA	inst460	(r13s[9], pp[217], r14c[7], r14s[8], r14c[8]);
FA	inst461	(r13s[10], pp[218], r14c[8], r14s[9], r14c[9]);
FA	inst462	(r13s[11], pp[219], r14c[9], r14s[10], r14c[10]);
FA	inst463	(r13s[12], pp[220], r14c[10], r14s[11], r14c[11]);
FA	inst464	(r13s[13], pp[221], r14c[11], r14s[12], r14c[12]);
FA	inst465	(r13s[14], pp[222], r14c[12], r14s[13], r14c[13]);
FA	inst466	(r13c[14], pp[223], r14c[13], r14s[14], r14c[14]);

HA	inst467	(r14s[1], pp[240], m[15], r15c[0]);
FA	inst468	(r14s[2], pp[226], r15c[0], r15s[1], r15c[1]);
FA	inst469	(r14s[3], pp[227], r15c[1], r15s[2], r15c[2]);
FA	inst470	(r14s[4], pp[228], r15c[2], r15s[3], r15c[3]);
FA	inst471	(r14s[5], pp[229], r15c[3], r15s[4], r15c[4]);
FA	inst472	(r14s[6], pp[230], r15c[4], r15s[5], r15c[5]);
FA	inst473	(r14s[7], pp[231], r15c[5], r15s[6], r15c[6]);
FA	inst474	(r14s[8], pp[232], r15c[6], r15s[7], r15c[7]);
FA	inst475	(r14s[9], pp[233], r15c[7], r15s[8], r15c[8]);
FA	inst476	(r14s[10], pp[234], r15c[8], r15s[9], r15c[9]);
FA	inst477	(r14s[11], pp[235], r15c[9], r15s[10], r15c[10]);
FA	inst478	(r14s[12], pp[236], r15c[10], r15s[11], r15c[11]);
FA	inst479	(r14s[13], pp[237], r15c[11], r15s[12], r15c[12]);
FA	inst480	(r14s[14], pp[238], r15c[12], r15s[13], r15c[13]);
FA	inst481	(r14c[14], pp[239], r15c[13], r15s[14], r15c[14]);

HA	inst482	(r15s[1], pp[241], m[16], r16c[0]);
FA	inst483	(r15s[2], pp[242], r16c[0], m[17], r16c[1]);
FA	inst484	(r15s[3], pp[243], r16c[1], m[18], r16c[2]);
FA	inst485	(r15s[4], pp[244], r16c[2], m[19], r16c[3]);
FA	inst486	(r15s[5], pp[245], r16c[3], m[20], r16c[4]);
FA	inst487	(r15s[6], pp[246], r16c[4], m[21], r16c[5]);
FA	inst488	(r15s[7], pp[247], r16c[5], m[22], r16c[6]);
FA	inst489	(r15s[8], pp[248], r16c[6], m[23], r16c[7]);
FA	inst490	(r15s[9], pp[249], r16c[7], m[24], r16c[8]);
FA	inst491	(r15s[10], pp[250], r16c[8], m[25], r16c[9]);
FA	inst492	(r15s[11], pp[251], r16c[9], m[26], r16c[10]);
FA	inst493	(r15s[12], pp[252], r16c[10], m[27], r16c[11]);
FA	inst494	(r15s[13], pp[253], r16c[11], m[28], r16c[12]);
FA	inst495	(r15s[14], pp[254], r16c[12], m[29], r16c[13]);
FA	inst496	(r15c[14], pp[255], r16c[13], m[30], m[31]);
endmodule

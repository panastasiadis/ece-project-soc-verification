VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 1000 ;
END UNITS

#USEMINSPACING OBS ON ;
#USEMINSPACING PIN OFF ;
#CLEARANCEMEASURE EUCLIDEAN ;


MANUFACTURINGGRID 0.005 ;

LAYER Metal1
  TYPE		ROUTING ;
  DIRECTION	HORIZONTAL ;
  PITCH		1.25  ;
  OFFSET	0  ;
  WIDTH		0.6 ;
  SPACING	0.5 ;
  RESISTANCE	RPERSQ 0.111 ;
  CAPACITANCE	CPERSQDIST 2.39e-05 ;
  EDGECAPACITANCE 0.0001776 ;
  HEIGHT 2.2 ;
  THICKNESS 0.63 ;
END Metal1

LAYER Via1
  TYPE	CUT ;
  SPACING	0.65 ;
END Via1

LAYER Metal2
  TYPE		ROUTING ;
  DIRECTION	VERTICAL ;
  PITCH		1.25  ;
  OFFSET	0  ;
  WIDTH		0.6 ;
  SPACING	0.65 ;
  RESISTANCE	RPERSQ 0.073 ;
  CAPACITANCE	CPERSQDIST 1.87e-05 ;
  EDGECAPACITANCE 0.000198 ;
  HEIGHT 3.73 ;
  THICKNESS 0.73 ;
END Metal2

LAYER Via2
  TYPE	CUT ;
  SPACING	0.65 ;
END Via2

LAYER Metal3
  TYPE		ROUTING ;
  DIRECTION	HORIZONTAL ;
  PITCH		1.25  ;
  WIDTH		0.6 ;
  SPACING	0.65 ;
  RESISTANCE	RPERSQ 0.078 ;
  CAPACITANCE	CPERSQDIST 1.5e-05 ;
  EDGECAPACITANCE 0.000197 ;
  HEIGHT 5.36 ;
  THICKNESS 0.705 ;
END Metal3

LAYER Via3
  TYPE	CUT ;
  SPACING	0.65 ;
END Via3

LAYER Metal4
  TYPE		ROUTING ;
  DIRECTION	VERTICAL ;
  PITCH		1.25  ;
  WIDTH		0.6 ;
  SPACING	0.65 ;
  RESISTANCE	RPERSQ 0.063 ;
  CAPACITANCE	CPERSQDIST 1.12e-05 ;
  EDGECAPACITANCE 0.000202 ;
  HEIGHT 6.97 ;
  THICKNESS 0.73 ;
END Metal4

LAYER Via4
  TYPE	CUT ;
  SPACING	0.65 ;
END Via4

LAYER Metal5
  TYPE		ROUTING ;
  DIRECTION	HORIZONTAL ;
  PITCH		1.25  ;
  WIDTH		0.6 ;
  SPACING	0.65 ;
  RESISTANCE	RPERSQ 0.063 ;
  CAPACITANCE	CPERSQDIST 1.11e-05 ;
  EDGECAPACITANCE 0.000202 ;
  HEIGHT 8.6 ;
  THICKNESS 0.73 ;
END Metal5

SPACING
  SAMENET Via1  Via1	0.65 ;
  SAMENET Via2  Via2	0.65 ;
  SAMENET Via3  Via3	0.65 ;
  SAMENET Via4  Via4	0.65 ;
  SAMENET Via1  Via2	0.00 ;
  SAMENET Via2  Via3	0.00 ;
  SAMENET Via3  Via4	0.00 ;
  SAMENET Metal2  Metal2	0.65 ;
  SAMENET Metal3  Metal3	0.65 ;
  SAMENET Metal4  Metal4	0.65 ;
  SAMENET Metal5  Metal5	0.65 ;
END SPACING

VIA ruleVia1 
  LAYER Metal1 ;
    RECT -0.400 -0.400 0.400 0.400 ;
  LAYER Via1 ;
    RECT -0.300 -0.300 0.300 0.300 ;
  LAYER Metal2 ;
    RECT -0.400 -0.400 0.400 0.400 ;
END ruleVia1

VIA ruleVia2 
  LAYER Metal2 ;
    RECT -0.300 -0.300 0.300 0.300 ;
  LAYER Via2 ;
    RECT -0.300 -0.300 0.300 0.300 ;
  LAYER Metal3 ;
    RECT -0.300 -0.300 0.300 0.300 ;
END ruleVia2

VIA ruleVia3 
  LAYER Metal3 ;
    RECT -0.300 -0.300 0.300 0.300 ;
  LAYER Via3 ;
    RECT -0.300 -0.300 0.300 0.300 ;
  LAYER Metal4 ;
    RECT -0.300 -0.300 0.300 0.300 ;
END ruleVia3

VIA ruleVia4 
  LAYER Metal4 ;
    RECT -0.300 -0.300 0.300 0.300 ;
  LAYER Via4 ;
    RECT -0.300 -0.300 0.300 0.300 ;
  LAYER Metal5 ;
    RECT -0.300 -0.300 0.300 0.300 ;
END ruleVia4

VIA M2_M1 DEFAULT
  LAYER Metal1 ;
    RECT -0.400 -0.400 0.400 0.400 ;
  LAYER Via1 ;
    RECT -0.300 -0.300 0.300 0.300 ;
  LAYER Metal2 ;
    RECT -0.300 -0.300 0.300 0.300 ;
  RESISTANCE 2.00 ;
END M2_M1

VIA M3_M2 DEFAULT
  LAYER Metal2 ;
    RECT -0.300 -0.300 0.300 0.300 ;
  LAYER Via2 ;
    RECT -0.300 -0.300 0.300 0.300 ;
  LAYER Metal3 ;
    RECT -0.300 -0.300 0.300 0.300 ;
  RESISTANCE 2.00 ;
END M3_M2

VIA M4_M3 DEFAULT
  LAYER Metal3 ;
    RECT -0.300 -0.300 0.300 0.300 ;
  LAYER Via3 ;
    RECT -0.300 -0.300 0.300 0.300 ;
  LAYER Metal4 ;
    RECT -0.300 -0.300 0.300 0.300 ;
  RESISTANCE 2.00 ;
END M4_M3

VIA M5_M4 DEFAULT
  LAYER Metal4 ;
    RECT -0.300 -0.300 0.300 0.300 ;
  LAYER Via4 ;
    RECT -0.300 -0.300 0.300 0.300 ;
  LAYER Metal5 ;
    RECT -0.300 -0.300 0.300 0.300 ;
  RESISTANCE 2.00 ;
END M5_M4

VIA M3_M2s DEFAULT
  TOPOFSTACKONLY
  LAYER Metal2 ;
    RECT -0.550 -0.550 0.550 0.550 ;
  LAYER Via2 ;
    RECT -0.300 -0.300 0.300 0.300 ;
  LAYER Metal3 ;
    RECT -0.300 -0.300 0.300 0.300 ;
  RESISTANCE 2.00 ;
END M3_M2s

VIA M4_M3s DEFAULT
  TOPOFSTACKONLY
  LAYER Metal3 ;
    RECT -0.550 -0.550 0.550 0.550 ;
  LAYER Via3 ;
    RECT -0.300 -0.300 0.300 0.300 ;
  LAYER Metal4 ;
    RECT -0.300 -0.300 0.300 0.300 ;
  RESISTANCE 2.00 ;
END M4_M3s

VIA M5_M4s DEFAULT
  TOPOFSTACKONLY
  LAYER Metal4 ;
    RECT -0.550 -0.550 0.550 0.550 ;
  LAYER Via4 ;
    RECT -0.300 -0.300 0.300 0.300 ;
  LAYER Metal5 ;
    RECT -0.300 -0.300 0.300 0.300 ;
  RESISTANCE 2.00 ;
END M5_M4s


VIARULE ruleVia1 GENERATE
  LAYER Metal1 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.1 ;
    METALOVERHANG 0 ;
  LAYER Metal2 ;
    DIRECTION VERTICAL ;
    OVERHANG 0 ;
    METALOVERHANG 0 ;
  LAYER Via1 ;
    RECT -0.3 -0.3 0.3 0.3 ;
    SPACING 1.25 BY 1.25 ;
END ruleVia1

VIARULE ruleVia2 GENERATE
  LAYER Metal2 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0 ;
    METALOVERHANG 0 ;
  LAYER Metal3 ;
    DIRECTION VERTICAL ;
    OVERHANG 0 ;
    METALOVERHANG 0 ;
  LAYER Via2 ;
    RECT -0.3 -0.3 0.3 0.3 ;
    SPACING 1.25 BY 1.25 ;
END ruleVia2

VIARULE ruleVia3 GENERATE
  LAYER Metal3 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0 ;
    METALOVERHANG 0 ;
  LAYER Metal4 ;
    DIRECTION VERTICAL ;
    OVERHANG 0 ;
    METALOVERHANG 0 ;
  LAYER Via3 ;
    RECT -0.3 -0.3 0.3 0.3 ;
    SPACING 1.25 BY 1.25 ;
    END ruleVia3

VIARULE ruleVia4 GENERATE
  LAYER Metal4 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0 ;
    METALOVERHANG 0 ;
  LAYER Metal5 ;
    DIRECTION VERTICAL ;
    OVERHANG 0 ;
    METALOVERHANG 0 ;
  LAYER Via4 ;
    RECT -0.3 -0.3 0.3 0.3 ;
    SPACING 1.25 BY 1.25 ;
END ruleVia4

VIARULE TURN1 GENERATE
  LAYER Metal1 ;
    DIRECTION HORIZONTAL ;
  LAYER Metal1 ;
    DIRECTION VERTICAL ;
END TURN1

VIARULE TURN2 GENERATE
  LAYER Metal2 ;
    DIRECTION HORIZONTAL ;
  LAYER Metal2 ;
    DIRECTION VERTICAL ;
END TURN2

VIARULE TURN3 GENERATE
  LAYER Metal3 ;
    DIRECTION HORIZONTAL ;
  LAYER Metal3 ;
    DIRECTION VERTICAL ;
END TURN3

VIARULE TURN4 GENERATE
  LAYER Metal4 ;
    DIRECTION HORIZONTAL ;
  LAYER Metal4 ;
    DIRECTION VERTICAL ;
END TURN4

VIARULE TURN5 GENERATE
  LAYER Metal5 ;
    DIRECTION HORIZONTAL ;
  LAYER Metal5 ;
    DIRECTION VERTICAL ;
END TURN5

SITE  core
    CLASS	CORE ;
    SYMMETRY	Y ;
    SIZE	1.250 BY 16.250 ;
END  core

SITE  io_site
    CLASS	PAD ;
    SYMMETRY	X ;
    SIZE	28.750 BY 600.000 ;
END  io_site

SITE  io_corner
    CLASS	PAD ;
    SYMMETRY	X Y ;
    SIZE	600.000 BY 600.000 ;
END  io_corner

SITE  CoreSite
    CLASS	CORE ;
    SYMMETRY	Y ;
    SIZE	1.250 BY 591.050 ;
END  CoreSite

MACRO tinvh_8
  CLASS  CORE ;
  FOREIGN tinvh_8 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 17.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.850 7.200 2.900 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 2.150 0.000 2.750 2.700 ;
        RECT 0.000 0.000 17.500 2.500 ;
        RECT 5.550 0.000 6.150 2.700 ;
    END
  END vss!
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 2.150 13.550 2.750 16.250 ;
        RECT 0.000 13.750 17.500 16.250 ;
        RECT 14.750 13.550 15.350 16.250 ;
        RECT 11.350 13.550 11.950 16.250 ;
    END
  END vdd!
  PIN en
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 14.200 7.200 16.550 7.800 ;
    END
  END en
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.950 7.200 10.400 7.800 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 3.800 5.950 6.350 6.550 ;
        RECT 8.850 5.950 13.650 6.550 ;
        RECT 13.050 5.950 13.650 7.800 ;
  END 
END tinvh_8

MACRO tinvh_7
  CLASS  CORE ;
  FOREIGN tinvh_7 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 16.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.850 7.200 2.900 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 2.150 0.000 2.750 2.700 ;
        RECT 0.000 0.000 16.250 2.500 ;
        RECT 9.500 0.000 10.100 2.700 ;
        RECT 5.850 0.000 6.450 2.700 ;
    END
  END vss!
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 2.150 13.550 2.750 16.250 ;
        RECT 0.000 13.750 16.250 16.250 ;
    END
  END vdd!
  PIN en
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 12.950 7.200 15.350 7.800 ;
    END
  END en
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.100 7.200 9.150 7.800 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 3.800 5.950 6.350 6.550 ;
        RECT 9.850 5.950 12.400 6.550 ;
        RECT 11.800 5.950 12.400 7.800 ;
  END 
END tinvh_7

MACRO tinvh_6
  CLASS  CORE ;
  FOREIGN tinvh_6 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.850 7.200 2.900 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 2.150 0.000 2.750 2.700 ;
        RECT 0.000 0.000 15.000 2.500 ;
    END
  END vss!
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 2.150 13.550 2.750 16.250 ;
        RECT 0.000 13.750 15.000 16.250 ;
    END
  END vdd!
  PIN en
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 11.700 7.200 14.100 7.800 ;
    END
  END en
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.200 7.200 8.200 7.800 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 3.800 5.900 6.350 6.550 ;
        RECT 8.650 5.950 11.150 6.550 ;
        RECT 10.550 5.950 11.150 7.800 ;
  END 
END tinvh_6

MACRO tinvh_5
  CLASS  CORE ;
  FOREIGN tinvh_5 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.850 7.200 2.900 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 2.150 0.000 2.750 2.700 ;
        RECT 0.000 0.000 15.000 2.500 ;
        RECT 5.550 0.000 6.150 2.700 ;
    END
  END vss!
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 2.150 13.550 2.750 16.250 ;
        RECT 0.000 13.750 15.000 16.250 ;
    END
  END vdd!
  PIN en
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 11.700 7.200 14.150 7.800 ;
    END
  END en
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.200 5.950 9.200 6.550 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 3.800 5.950 6.400 6.550 ;
        RECT 8.650 7.200 11.200 7.800 ;
  END 
END tinvh_5

MACRO tinvh_4
  CLASS  CORE ;
  FOREIGN tinvh_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.850 7.200 2.850 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 2.150 0.000 2.750 2.700 ;
        RECT 0.000 0.000 15.000 2.500 ;
        RECT 5.550 0.000 6.150 2.700 ;
    END
  END vss!
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 2.150 13.550 2.750 16.250 ;
        RECT 0.000 13.750 15.000 16.250 ;
    END
  END vdd!
  PIN en
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 11.700 7.200 14.150 7.800 ;
    END
  END en
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.200 5.950 9.200 6.550 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 3.800 5.950 6.300 6.550 ;
        RECT 8.650 7.200 11.200 7.800 ;
  END 
END tinvh_4

MACRO tinvh_3
  CLASS  CORE ;
  FOREIGN tinvh_3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.850 7.200 2.900 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 2.150 0.000 2.750 2.700 ;
        RECT 0.000 0.000 13.750 2.500 ;
        RECT 5.400 0.000 6.000 2.650 ;
    END
  END vss!
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 2.150 13.550 2.750 16.250 ;
        RECT 0.000 13.750 13.750 16.250 ;
    END
  END vdd!
  PIN en
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 10.250 7.200 12.800 7.800 ;
    END
  END en
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.950 5.950 6.550 9.100 ;
        RECT 5.950 5.950 7.800 6.550 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 3.800 5.950 5.350 6.550 ;
        RECT 4.700 5.950 5.350 9.100 ;
        RECT 7.150 7.200 9.000 7.800 ;
        RECT 8.400 5.950 9.000 9.050 ;
        RECT 8.400 8.450 9.900 9.050 ;
  END 
END tinvh_3

MACRO tinvh_2
  CLASS  CORE ;
  FOREIGN tinvh_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.850 7.200 2.850 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 2.150 0.000 2.750 2.700 ;
        RECT 0.000 0.000 13.750 2.500 ;
    END
  END vss!
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 2.150 13.550 2.750 16.250 ;
        RECT 0.000 13.750 13.750 16.250 ;
    END
  END vdd!
  PIN en
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 10.250 7.200 12.800 7.800 ;
    END
  END en
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.050 7.100 6.650 9.050 ;
        RECT 6.050 7.100 7.800 7.900 ;
        RECT 7.100 5.900 7.800 7.900 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 3.800 5.900 6.550 6.600 ;
        RECT 4.750 5.900 5.350 9.050 ;
        RECT 8.400 5.900 9.000 9.050 ;
        RECT 7.150 8.400 9.950 9.050 ;
  END 
END tinvh_2

MACRO tinvh_16
  CLASS  CORE ;
  FOREIGN tinvh_16 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 20.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.850 7.200 2.900 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 2.150 0.000 2.750 2.700 ;
        RECT 0.000 0.000 20.000 2.500 ;
        RECT 8.950 0.000 9.550 2.650 ;
        RECT 5.550 0.000 6.150 2.700 ;
    END
  END vss!
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 2.100 13.550 2.800 16.250 ;
        RECT 0.000 13.750 20.000 16.250 ;
        RECT 14.100 13.550 14.800 16.250 ;
        RECT 10.700 13.550 11.400 16.250 ;
        RECT 7.300 13.550 8.000 16.250 ;
    END
  END vdd!
  PIN en
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 16.700 7.200 19.050 7.800 ;
    END
  END en
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.000 8.450 13.100 9.050 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 3.750 5.950 6.600 6.550 ;
        RECT 3.750 5.950 4.350 9.100 ;
        RECT 3.750 8.400 5.350 9.100 ;
        RECT 13.700 5.900 15.450 6.600 ;
        RECT 14.800 5.900 15.450 7.900 ;
        RECT 14.800 7.200 16.200 7.900 ;
        RECT 4.850 7.150 14.300 7.850 ;
        RECT 13.600 7.150 14.300 9.050 ;
        RECT 13.600 8.450 19.550 9.050 ;
  END 
END tinvh_16

MACRO tinvh_14
  CLASS  CORE ;
  FOREIGN tinvh_14 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 18.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.850 7.200 2.900 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 2.150 0.000 2.750 2.700 ;
        RECT 0.000 0.000 18.750 2.500 ;
        RECT 5.550 0.000 6.150 2.700 ;
    END
  END vss!
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 2.150 13.550 2.750 16.250 ;
        RECT 0.000 13.750 18.750 16.250 ;
        RECT 12.600 13.550 13.200 16.250 ;
        RECT 9.200 13.550 9.800 16.250 ;
    END
  END vdd!
  PIN en
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 15.450 7.200 17.800 7.800 ;
    END
  END en
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.450 8.450 11.550 9.050 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 3.500 5.900 6.350 6.600 ;
        RECT 3.500 5.900 4.100 9.100 ;
        RECT 3.500 8.400 5.400 9.100 ;
        RECT 12.550 5.950 14.900 6.550 ;
        RECT 14.300 5.950 14.900 8.000 ;
        RECT 4.600 7.150 13.700 7.850 ;
        RECT 13.000 7.150 13.700 9.100 ;
        RECT 17.650 8.400 18.350 9.100 ;
        RECT 13.000 8.500 18.350 9.100 ;
  END 
END tinvh_14

MACRO tinvh_12
  CLASS  CORE ;
  FOREIGN tinvh_12 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 18.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.850 7.200 2.900 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 2.150 0.000 2.750 2.700 ;
        RECT 0.000 0.000 18.750 2.500 ;
        RECT 9.200 0.000 9.800 2.650 ;
        RECT 5.700 0.000 6.300 2.700 ;
    END
  END vss!
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 2.150 13.550 2.750 16.250 ;
        RECT 0.000 13.750 18.750 16.250 ;
        RECT 12.600 13.550 13.200 16.250 ;
        RECT 9.200 13.550 9.800 16.250 ;
    END
  END vdd!
  PIN en
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 15.450 7.200 17.900 7.800 ;
    END
  END en
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.450 8.450 11.650 9.050 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 3.800 5.900 10.450 6.500 ;
        RECT 3.800 5.900 4.500 9.050 ;
        RECT 3.800 8.450 5.350 9.050 ;
        RECT 12.550 5.900 14.950 6.600 ;
        RECT 14.250 5.900 14.950 7.950 ;
        RECT 5.100 7.250 13.600 7.850 ;
        RECT 13.000 7.250 13.600 9.050 ;
        RECT 13.000 8.450 18.350 9.050 ;
  END 
END tinvh_12

MACRO tinvh_10
  CLASS  CORE ;
  FOREIGN tinvh_10 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 17.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.850 7.200 2.850 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 2.150 0.000 2.750 2.700 ;
        RECT 0.000 0.000 17.500 2.500 ;
        RECT 8.950 0.000 9.550 2.650 ;
        RECT 5.550 0.000 6.150 2.700 ;
    END
  END vss!
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 2.150 13.550 2.750 16.250 ;
        RECT 0.000 13.750 17.500 16.250 ;
        RECT 11.350 13.550 11.950 16.250 ;
        RECT 7.950 13.550 8.550 16.250 ;
    END
  END vdd!
  PIN en
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 14.200 7.200 16.650 7.800 ;
    END
  END en
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.200 8.450 10.300 9.050 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 3.850 6.150 4.450 9.050 ;
        RECT 3.850 8.450 5.350 9.050 ;
        RECT 8.350 5.900 13.700 6.600 ;
        RECT 13.000 5.900 13.700 7.950 ;
        RECT 5.100 7.000 5.800 7.850 ;
        RECT 5.100 7.150 12.350 7.850 ;
        RECT 11.750 7.150 12.350 9.050 ;
        RECT 11.750 8.450 17.100 9.050 ;
  END 
END tinvh_10

MACRO tinvh_1
  CLASS  CORE ;
  FOREIGN tinvh_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 8.450 2.250 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 11.250 2.500 ;
    END
  END vss!
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 1.000 13.550 1.600 16.250 ;
        RECT 0.000 13.750 11.250 16.250 ;
    END
  END vdd!
  PIN en
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.750 7.200 10.750 7.800 ;
    END
  END en
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.900 5.950 5.500 9.150 ;
        RECT 4.900 5.950 6.750 6.550 ;
        RECT 4.900 5.950 5.850 6.650 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 2.700 5.850 4.350 6.450 ;
        RECT 3.750 5.850 4.350 8.350 ;
        RECT 2.700 3.400 7.850 4.050 ;
        RECT 7.350 5.900 8.050 9.100 ;
        RECT 6.200 8.500 8.900 9.100 ;
  END 
END tinvh_1

MACRO tbufh_8
  CLASS  CORE ;
  FOREIGN tbufh_8 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 18.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.550 7.200 2.600 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 18.750 2.500 ;
    END
  END vss!
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 8.950 13.550 9.550 16.250 ;
        RECT 0.000 13.750 18.750 16.250 ;
        RECT 12.350 13.550 12.950 16.250 ;
    END
  END vdd!
  PIN en
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 15.200 7.200 17.200 7.800 ;
    END
  END en
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.250 7.200 11.300 7.800 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 2.400 5.900 6.700 6.600 ;
        RECT 3.350 5.900 3.950 9.050 ;
        RECT 11.900 7.200 14.700 7.800 ;
        RECT 4.600 7.150 5.300 9.100 ;
        RECT 4.600 8.400 18.100 9.100 ;
  END 
END tbufh_8

MACRO tbufh_7
  CLASS  CORE ;
  FOREIGN tbufh_7 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.300 7.200 2.300 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 3.850 0.000 4.450 2.700 ;
        RECT 0.000 0.000 15.000 2.500 ;
    END
  END vss!
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 15.000 16.250 ;
    END
  END vdd!
  PIN en
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 11.700 7.200 13.700 7.800 ;
    END
  END en
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.550 4.700 6.150 6.550 ;
        RECT 5.550 5.950 8.000 6.550 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 2.100 5.900 5.000 6.600 ;
        RECT 3.000 5.900 3.600 9.050 ;
        RECT 3.000 8.450 3.650 9.050 ;
        RECT 8.600 5.900 11.200 6.600 ;
        RECT 10.500 5.900 11.200 7.850 ;
        RECT 4.300 7.150 8.150 7.850 ;
        RECT 7.450 7.150 8.150 9.100 ;
        RECT 7.450 8.400 14.600 9.100 ;
  END 
END tbufh_7

MACRO tbufh_6
  CLASS  CORE ;
  FOREIGN tbufh_6 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.300 7.200 2.300 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 3.850 0.000 4.450 2.700 ;
        RECT 0.000 0.000 15.000 2.500 ;
    END
  END vss!
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 15.000 16.250 ;
    END
  END vdd!
  PIN en
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 11.700 7.200 13.700 7.800 ;
    END
  END en
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.500 5.950 8.000 6.550 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 2.100 5.950 5.000 6.550 ;
        RECT 3.050 5.950 3.650 9.050 ;
        RECT 8.650 7.200 11.200 7.800 ;
        RECT 4.350 7.250 8.150 7.850 ;
        RECT 7.450 7.250 8.150 9.100 ;
        RECT 7.450 8.450 14.600 9.100 ;
  END 
END tbufh_6

MACRO tbufh_5
  CLASS  CORE ;
  FOREIGN tbufh_5 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.300 7.200 2.300 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 3.850 0.000 4.450 2.700 ;
        RECT 0.000 0.000 13.750 2.500 ;
    END
  END vss!
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 4.350 13.550 4.950 16.250 ;
        RECT 0.000 13.750 13.750 16.250 ;
    END
  END vdd!
  PIN en
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 10.450 7.200 12.450 7.800 ;
    END
  END en
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.500 5.950 7.500 6.550 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 2.100 5.900 5.000 6.600 ;
        RECT 4.300 5.900 5.000 6.850 ;
        RECT 7.400 7.200 9.950 7.800 ;
  END 
END tbufh_5

MACRO tbufh_4
  CLASS  CORE ;
  FOREIGN tbufh_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.300 7.200 2.300 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 3.850 0.000 4.450 2.700 ;
        RECT 0.000 0.000 13.750 2.500 ;
    END
  END vss!
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 4.350 13.550 4.950 16.250 ;
        RECT 0.000 13.750 13.750 16.250 ;
    END
  END vdd!
  PIN en
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 10.450 7.200 12.450 7.800 ;
    END
  END en
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.500 5.950 7.500 6.550 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 2.100 5.900 5.000 6.600 ;
        RECT 7.400 7.200 9.950 7.800 ;
  END 
END tbufh_4

MACRO tbufh_3
  CLASS  CORE ;
  FOREIGN tbufh_3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.450 7.200 2.450 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 4.000 0.000 4.600 2.650 ;
        RECT 0.000 0.000 12.500 2.500 ;
    END
  END vss!
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 12.500 16.250 ;
    END
  END vdd!
  PIN en
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.850 7.200 10.850 7.800 ;
    END
  END en
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.450 5.950 5.150 9.100 ;
        RECT 4.450 5.950 6.350 6.550 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 2.250 5.900 3.850 6.600 ;
        RECT 3.150 5.900 3.850 9.100 ;
        RECT 5.650 7.150 7.650 7.850 ;
        RECT 6.950 5.900 7.650 9.100 ;
        RECT 6.950 8.400 8.550 9.100 ;
  END 
END tbufh_3

MACRO tbufh_16
  CLASS  CORE ;
  FOREIGN tbufh_16 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 21.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 7.200 2.300 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 8.550 0.000 9.150 2.650 ;
        RECT 0.000 0.000 21.250 2.500 ;
    END
  END vss!
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 8.300 13.550 8.900 16.250 ;
        RECT 0.000 13.750 21.250 16.250 ;
        RECT 15.100 13.550 15.700 16.250 ;
        RECT 11.700 13.550 12.300 16.250 ;
    END
  END vdd!
  PIN en
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 17.950 7.200 19.950 7.800 ;
    END
  END en
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.100 5.950 14.150 6.550 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 2.100 5.950 6.100 6.550 ;
        RECT 3.050 5.950 3.650 9.050 ;
        RECT 14.650 7.250 17.450 7.850 ;
        RECT 4.350 7.150 4.950 9.050 ;
        RECT 4.350 8.450 20.850 9.050 ;
  END 
END tbufh_16

MACRO tbufh_14
  CLASS  CORE ;
  FOREIGN tbufh_14 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 18.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.400 7.200 2.450 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 8.700 0.000 9.300 2.650 ;
        RECT 0.000 0.000 18.750 2.500 ;
    END
  END vss!
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 9.200 13.550 9.800 16.250 ;
        RECT 0.000 13.750 18.750 16.250 ;
        RECT 12.600 13.550 13.200 16.250 ;
    END
  END vdd!
  PIN en
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 15.450 7.200 17.450 7.800 ;
    END
  END en
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.500 5.950 11.500 6.550 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 2.000 5.900 6.550 6.600 ;
        RECT 3.200 5.900 3.800 9.050 ;
        RECT 12.150 7.200 14.950 7.800 ;
        RECT 4.500 7.150 5.100 9.050 ;
        RECT 4.500 8.450 18.350 9.050 ;
  END 
END tbufh_14

MACRO tbufh_12
  CLASS  CORE ;
  FOREIGN tbufh_12 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 18.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.400 7.200 2.450 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 9.200 0.000 9.800 2.650 ;
        RECT 0.000 0.000 18.750 2.500 ;
    END
  END vss!
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 9.200 13.550 9.800 16.250 ;
        RECT 0.000 13.750 18.750 16.250 ;
        RECT 12.600 13.550 13.200 16.250 ;
    END
  END vdd!
  PIN en
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 15.450 7.200 17.450 7.800 ;
    END
  END en
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.500 7.200 11.550 7.800 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 2.000 5.900 10.450 6.600 ;
        RECT 3.200 5.900 3.800 9.050 ;
        RECT 12.150 7.150 14.950 7.800 ;
        RECT 4.450 7.150 5.050 9.100 ;
        RECT 4.450 8.400 18.350 9.100 ;
  END 
END tbufh_12

MACRO tbufh_10
  CLASS  CORE ;
  FOREIGN tbufh_10 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 18.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.550 7.200 2.600 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 8.950 0.000 9.550 2.650 ;
        RECT 0.000 0.000 18.750 2.500 ;
    END
  END vss!
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 8.950 13.550 9.550 16.250 ;
        RECT 0.000 13.750 18.750 16.250 ;
        RECT 12.350 13.550 12.950 16.250 ;
    END
  END vdd!
  PIN en
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 15.200 7.200 17.200 7.800 ;
    END
  END en
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.100 5.950 11.300 6.550 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 2.000 5.950 6.600 6.550 ;
        RECT 3.350 5.950 3.950 9.050 ;
        RECT 11.900 7.150 14.700 7.800 ;
        RECT 4.600 7.150 5.300 9.100 ;
        RECT 4.600 8.400 18.100 9.100 ;
  END 
END tbufh_10

MACRO tbufh_2
  CLASS  CORE ;
  FOREIGN tbufh_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 8.450 2.250 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 3.750 0.000 4.350 2.700 ;
        RECT 0.000 0.000 10.000 2.500 ;
    END
  END vss!
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 5.950 13.550 6.550 16.250 ;
        RECT 0.000 13.750 10.000 16.250 ;
    END
  END vdd!
  PIN en
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.750 7.200 9.750 7.800 ;
    END
  END en
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.250 5.950 4.850 9.150 ;
        RECT 4.250 5.950 5.750 6.550 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 2.000 5.800 2.700 7.850 ;
        RECT 2.000 7.150 3.750 7.850 ;
        RECT 3.050 7.150 3.750 8.400 ;
        RECT 1.900 3.400 6.850 4.100 ;
        RECT 6.350 5.900 7.050 9.150 ;
        RECT 5.350 8.450 7.950 9.150 ;
  END 
END tbufh_2

MACRO tbufh_1
  CLASS  CORE ;
  FOREIGN tbufh_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 8.450 2.250 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 10.000 2.500 ;
    END
  END vss!
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 10.000 16.250 ;
    END
  END vdd!
  PIN en
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.750 7.200 9.750 7.800 ;
    END
  END en
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.250 5.950 4.850 9.150 ;
        RECT 4.250 5.950 5.750 6.550 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 2.000 5.800 2.700 7.850 ;
        RECT 2.000 7.150 3.750 7.850 ;
        RECT 3.050 7.150 3.750 8.400 ;
        RECT 1.900 3.400 6.850 4.100 ;
        RECT 6.350 5.900 7.050 9.150 ;
        RECT 5.400 8.450 7.950 9.150 ;
  END 
END tbufh_1

MACRO sdffpt_8
  CLASS  CORE ;
  FOREIGN sdffpt_8 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 36.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 30.750 5.950 32.750 6.550 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 36.250 2.500 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.350 7.200 7.150 7.800 ;
    END
  END d
  PIN se
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.350 8.450 4.850 9.050 ;
    END
  END se
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 1.000 13.450 1.600 16.250 ;
        RECT 0.000 13.750 36.250 16.250 ;
        RECT 26.500 13.450 27.100 16.250 ;
        RECT 8.400 13.450 9.000 16.250 ;
    END
  END vdd!
  PIN setb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.100 5.950 3.100 6.550 ;
    END
  END setb
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 26.800 8.450 29.300 9.050 ;
    END
  END qb
  PIN sdi
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.750 4.700 11.750 5.300 ;
    END
  END sdi
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 33.700 4.700 35.750 5.300 ;
    END
  END ck
  OBS 
      LAYER Metal1 ;
        RECT 3.950 6.000 8.250 6.600 ;
        RECT 7.650 6.000 8.250 7.950 ;
        RECT 7.650 7.350 10.300 7.950 ;
        RECT 2.150 9.700 12.100 10.300 ;
        RECT 13.200 5.500 13.800 10.300 ;
        RECT 13.200 9.700 14.900 10.300 ;
        RECT 14.400 5.950 21.850 6.550 ;
        RECT 14.400 5.950 15.000 8.950 ;
        RECT 14.400 8.350 19.200 8.950 ;
        RECT 17.300 9.500 25.400 10.100 ;
        RECT 19.700 4.700 30.900 5.300 ;
        RECT 15.500 7.250 35.600 7.850 ;
  END 
END sdffpt_8

MACRO sdffpt_6
  CLASS  CORE ;
  FOREIGN sdffpt_6 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 35.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 29.500 9.700 31.500 10.300 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 28.800 0.000 29.400 2.650 ;
        RECT 0.000 0.000 35.000 2.500 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.000 7.200 6.600 7.800 ;
    END
  END d
  PIN se
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.400 8.450 4.100 9.050 ;
    END
  END se
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 1.000 13.450 1.600 16.250 ;
        RECT 0.000 13.750 35.000 16.250 ;
        RECT 28.800 13.450 29.400 16.250 ;
        RECT 7.750 13.450 8.350 16.250 ;
    END
  END vdd!
  PIN setb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.900 5.950 2.900 6.550 ;
    END
  END setb
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 24.100 8.450 26.100 9.050 ;
    END
  END qb
  PIN sdi
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.400 4.650 11.100 5.450 ;
    END
  END sdi
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 32.500 5.950 34.500 6.550 ;
    END
  END ck
  OBS 
      LAYER Metal1 ;
        RECT 3.450 6.000 7.750 6.600 ;
        RECT 7.150 6.000 7.750 7.800 ;
        RECT 7.150 7.200 9.250 7.800 ;
        RECT 2.850 4.750 8.850 5.350 ;
        RECT 8.250 4.750 8.850 6.650 ;
        RECT 8.250 6.050 11.200 6.650 ;
        RECT 10.000 6.050 10.600 10.300 ;
        RECT 2.750 9.700 11.300 10.300 ;
        RECT 11.800 4.900 12.900 5.500 ;
        RECT 11.800 4.900 12.400 10.350 ;
        RECT 11.800 9.750 14.000 10.350 ;
        RECT 20.100 5.950 20.700 6.700 ;
        RECT 13.150 6.100 20.700 6.700 ;
        RECT 13.150 6.100 13.750 9.250 ;
        RECT 13.150 8.600 18.100 9.200 ;
        RECT 13.150 8.600 14.350 9.250 ;
        RECT 18.800 9.650 27.700 10.250 ;
        RECT 16.200 9.700 19.400 10.300 ;
        RECT 22.750 7.100 29.000 7.700 ;
        RECT 22.750 7.100 23.350 9.150 ;
        RECT 18.600 8.550 23.350 9.150 ;
        RECT 21.650 6.000 30.750 6.600 ;
        RECT 30.150 6.000 30.750 7.800 ;
        RECT 14.250 7.200 22.250 7.800 ;
        RECT 30.150 7.200 34.550 7.800 ;
        RECT 21.650 6.000 22.250 7.850 ;
        RECT 19.700 7.200 22.250 7.850 ;
        RECT 14.250 7.200 14.850 8.000 ;
  END 
END sdffpt_6

MACRO sdffpt_4
  CLASS  CORE ;
  FOREIGN sdffpt_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 32.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 28.050 7.200 30.050 7.800 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 32.500 2.500 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.000 8.200 4.600 9.050 ;
        RECT 2.600 8.450 4.600 9.050 ;
    END
  END d
  PIN se
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.850 4.700 6.850 5.300 ;
    END
  END se
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 2.150 13.550 2.750 16.250 ;
        RECT 0.000 13.750 32.500 16.250 ;
        RECT 15.300 13.550 15.900 16.250 ;
    END
  END vdd!
  PIN setb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.300 7.200 2.450 7.800 ;
    END
  END setb
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 24.250 5.950 26.250 6.550 ;
    END
  END qb
  PIN sdi
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.800 4.700 9.850 5.300 ;
    END
  END sdi
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 15.050 5.950 17.000 6.550 ;
        RECT 16.400 5.950 17.000 6.950 ;
    END
  END ck
  OBS 
      LAYER Metal1 ;
        RECT 6.450 6.000 7.050 6.750 ;
        RECT 3.500 6.150 7.050 6.750 ;
        RECT 5.100 6.150 5.700 10.150 ;
        RECT 8.150 7.250 10.600 7.850 ;
        RECT 8.150 6.000 8.750 8.900 ;
        RECT 6.800 8.300 8.750 8.900 ;
        RECT 11.100 6.000 13.300 6.600 ;
        RECT 11.100 6.000 11.700 10.150 ;
        RECT 11.100 9.550 13.100 10.150 ;
        RECT 18.050 6.350 23.600 6.950 ;
        RECT 13.200 7.250 15.900 7.850 ;
        RECT 18.050 6.300 18.650 8.050 ;
        RECT 15.300 7.450 18.650 8.050 ;
        RECT 12.200 8.350 12.800 9.050 ;
        RECT 12.200 8.450 14.800 9.050 ;
        RECT 19.700 8.450 24.250 9.050 ;
        RECT 19.700 7.950 20.300 9.150 ;
        RECT 14.200 8.550 20.300 9.150 ;
  END 
END sdffpt_4

MACRO sdffpt_3
  CLASS  CORE ;
  FOREIGN sdffpt_3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 28.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 24.800 5.950 26.800 6.550 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.950 0.000 1.650 2.700 ;
        RECT 0.000 0.000 28.750 2.500 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.300 8.450 4.300 9.050 ;
    END
  END d
  PIN se
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.550 4.650 6.550 5.300 ;
    END
  END se
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 1.850 13.550 2.450 16.250 ;
        RECT 0.000 13.750 28.750 16.250 ;
    END
  END vdd!
  PIN setb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.300 7.200 2.300 7.800 ;
    END
  END setb
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 22.000 5.950 24.000 6.550 ;
    END
  END qb
  PIN sdi
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.250 4.700 9.250 5.300 ;
    END
  END sdi
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 15.200 5.950 17.200 6.550 ;
    END
  END ck
  OBS 
      LAYER Metal1 ;
        RECT 3.100 6.000 6.300 6.600 ;
        RECT 4.800 6.000 5.400 9.300 ;
        RECT 7.400 7.250 9.700 7.850 ;
        RECT 7.400 6.000 8.000 9.200 ;
        RECT 6.500 8.600 8.000 9.200 ;
        RECT 10.200 5.950 12.050 6.550 ;
        RECT 10.200 5.950 10.800 10.150 ;
        RECT 10.200 9.550 12.100 10.150 ;
        RECT 11.300 8.450 21.700 9.050 ;
        RECT 12.100 7.350 21.700 7.950 ;
  END 
END sdffpt_3

MACRO sdffpt_2
  CLASS  CORE ;
  FOREIGN sdffpt_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 26.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 21.050 8.450 23.050 9.050 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 14.050 0.000 14.650 2.700 ;
        RECT 0.000 0.000 26.250 2.500 ;
        RECT 20.050 0.000 20.650 2.800 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.050 5.950 4.050 6.550 ;
        RECT 3.450 5.950 4.050 6.800 ;
    END
  END d
  PIN se
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.700 3.200 6.150 4.050 ;
    END
  END se
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 1.000 13.550 1.600 16.250 ;
        RECT 0.000 13.750 26.250 16.250 ;
        RECT 14.150 13.550 14.750 16.250 ;
    END
  END vdd!
  PIN setb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 8.450 2.250 9.050 ;
    END
  END setb
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 18.200 8.450 20.200 9.050 ;
    END
  END qb
  PIN sdi
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.050 8.400 8.950 9.100 ;
    END
  END sdi
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 23.750 8.450 25.750 9.050 ;
    END
  END ck
  OBS 
      LAYER Metal1 ;
        RECT 4.700 5.800 5.850 6.400 ;
        RECT 4.700 5.800 5.300 7.900 ;
        RECT 2.150 7.300 5.300 7.900 ;
        RECT 3.900 7.300 4.500 9.200 ;
        RECT 8.350 5.300 9.300 5.900 ;
        RECT 8.350 5.300 8.950 7.500 ;
        RECT 5.800 6.900 8.950 7.500 ;
        RECT 5.800 6.900 6.400 9.200 ;
        RECT 5.600 8.600 6.400 9.200 ;
        RECT 10.350 5.800 11.000 6.400 ;
        RECT 9.450 6.400 10.950 7.000 ;
        RECT 9.450 6.400 10.050 9.200 ;
        RECT 9.450 8.600 11.850 9.200 ;
        RECT 12.250 6.250 16.350 6.850 ;
        RECT 11.450 6.900 12.850 7.500 ;
        RECT 12.250 6.250 12.850 7.500 ;
        RECT 10.550 7.500 12.050 8.100 ;
        RECT 17.050 7.250 25.850 7.850 ;
        RECT 14.450 7.350 17.650 7.950 ;
        RECT 14.450 7.350 15.050 8.600 ;
        RECT 12.550 8.000 15.050 8.600 ;
  END 
END sdffpt_2

MACRO sdffpt_1
  CLASS  CORE ;
  FOREIGN sdffpt_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 25.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 22.750 5.950 24.750 6.550 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 16.200 0.000 16.800 2.700 ;
        RECT 0.000 0.000 25.000 2.500 ;
        RECT 22.350 0.000 22.950 2.700 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.150 5.900 4.050 6.800 ;
    END
  END d
  PIN se
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.600 3.200 6.150 4.050 ;
    END
  END se
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 1.000 13.550 1.600 16.250 ;
        RECT 0.000 13.750 25.000 16.250 ;
        RECT 22.250 13.550 22.850 16.250 ;
        RECT 14.450 13.550 15.050 16.250 ;
    END
  END vdd!
  PIN setb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 8.450 2.250 9.050 ;
    END
  END setb
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 22.000 8.450 24.000 9.050 ;
    END
  END qb
  PIN sdi
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.900 8.350 8.400 9.150 ;
    END
  END sdi
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 14.050 3.450 16.050 4.050 ;
    END
  END ck
  OBS 
      LAYER Metal1 ;
        RECT 4.550 5.800 5.850 6.400 ;
        RECT 4.550 5.800 5.150 7.900 ;
        RECT 2.150 7.300 5.150 7.900 ;
        RECT 3.900 7.300 4.500 9.200 ;
        RECT 7.800 5.300 9.300 5.900 ;
        RECT 7.800 5.300 8.400 7.500 ;
        RECT 5.650 6.900 8.400 7.500 ;
        RECT 5.650 6.900 6.250 9.200 ;
        RECT 5.600 8.600 6.250 9.200 ;
        RECT 9.800 5.800 11.100 6.400 ;
        RECT 8.900 6.400 10.400 7.000 ;
        RECT 8.900 6.400 9.500 9.200 ;
        RECT 8.900 8.600 11.900 9.200 ;
        RECT 11.750 6.250 17.800 6.850 ;
        RECT 11.100 6.950 12.350 7.550 ;
        RECT 11.750 6.250 12.350 7.550 ;
        RECT 10.000 7.500 11.700 8.100 ;
        RECT 17.200 8.450 20.400 9.050 ;
        RECT 15.900 7.350 21.100 7.950 ;
        RECT 15.900 7.350 16.500 8.950 ;
        RECT 12.450 8.350 16.500 8.950 ;
  END 
END sdffpt_1

MACRO sdffps_8
  CLASS  CORE ;
  FOREIGN sdffps_8 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 35.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN sb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.300 7.150 1.800 7.950 ;
    END
  END sb
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 23.450 8.450 27.950 9.050 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 20.450 0.000 21.050 2.800 ;
        RECT 0.000 0.000 35.000 2.500 ;
        RECT 25.150 0.000 25.750 2.800 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.400 5.950 5.350 6.550 ;
        RECT 4.750 5.950 5.350 6.700 ;
    END
  END d
  PIN se
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.200 8.450 2.800 9.150 ;
        RECT 2.200 8.450 7.450 9.050 ;
    END
  END se
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 5.700 13.450 6.300 16.250 ;
        RECT 0.000 13.750 35.000 16.250 ;
        RECT 25.150 13.450 25.750 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 29.400 9.700 31.400 10.300 ;
    END
  END qb
  PIN sdi
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.200 4.700 8.700 5.650 ;
    END
  END sdi
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 32.350 4.700 34.350 5.300 ;
    END
  END ck
  OBS 
      LAYER Metal1 ;
        RECT 2.350 7.250 6.150 7.850 ;
        RECT 1.950 4.550 6.550 5.150 ;
        RECT 5.950 4.550 6.550 6.750 ;
        RECT 5.950 6.150 9.450 6.750 ;
        RECT 8.850 6.150 9.450 10.300 ;
        RECT 1.600 9.700 9.450 10.300 ;
        RECT 9.950 5.000 11.150 5.600 ;
        RECT 9.950 5.000 10.550 10.300 ;
        RECT 9.950 9.700 11.200 10.300 ;
        RECT 12.650 6.050 19.100 6.650 ;
        RECT 11.250 6.100 13.250 6.750 ;
        RECT 11.250 6.100 11.850 9.150 ;
        RECT 13.450 8.450 16.150 9.050 ;
        RECT 11.050 8.550 14.050 9.150 ;
        RECT 14.250 9.650 22.750 10.250 ;
        RECT 16.650 4.700 25.300 5.300 ;
        RECT 28.950 5.700 29.550 6.550 ;
        RECT 23.400 5.950 29.550 6.550 ;
        RECT 20.500 7.200 34.250 7.800 ;
        RECT 12.350 7.350 21.100 7.950 ;
        RECT 12.350 7.350 12.950 8.050 ;
  END 
END sdffps_8

MACRO sdffps_6
  CLASS  CORE ;
  FOREIGN sdffps_6 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 32.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN sb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.950 8.850 1.550 10.300 ;
        RECT 0.350 9.700 1.550 10.300 ;
    END
  END sb
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 27.350 9.700 29.350 10.300 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 20.250 0.000 20.850 2.800 ;
        RECT 0.000 0.000 32.500 2.500 ;
        RECT 23.650 0.000 24.250 2.800 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.300 5.950 5.350 6.550 ;
    END
  END d
  PIN se
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.050 7.250 7.650 9.050 ;
        RECT 2.750 8.450 7.650 9.050 ;
    END
  END se
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 5.800 13.450 6.400 16.250 ;
        RECT 0.000 13.750 32.500 16.250 ;
        RECT 26.650 13.450 27.250 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 20.550 5.950 22.550 6.550 ;
    END
  END qb
  PIN sdi
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.000 4.700 9.000 5.300 ;
    END
  END sdi
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 30.100 8.450 32.100 9.050 ;
    END
  END ck
  OBS 
      LAYER Metal1 ;
        RECT 2.250 7.250 6.550 7.850 ;
        RECT 5.950 7.250 6.550 7.950 ;
        RECT 1.850 4.550 6.450 5.150 ;
        RECT 5.850 4.550 6.450 6.750 ;
        RECT 5.850 6.150 9.150 6.750 ;
        RECT 8.550 6.150 9.150 10.300 ;
        RECT 2.250 9.700 9.350 10.300 ;
        RECT 9.850 4.700 11.150 5.300 ;
        RECT 9.850 4.700 10.450 10.300 ;
        RECT 9.850 9.700 11.250 10.300 ;
        RECT 18.450 5.850 19.050 6.650 ;
        RECT 10.950 6.050 19.050 6.650 ;
        RECT 10.950 6.050 11.550 9.200 ;
        RECT 13.150 8.250 15.950 8.850 ;
        RECT 10.950 8.600 13.750 9.200 ;
        RECT 14.250 9.350 14.850 10.250 ;
        RECT 14.250 9.650 25.550 10.250 ;
        RECT 23.850 4.700 27.300 5.300 ;
        RECT 23.850 4.700 24.450 6.550 ;
        RECT 16.450 8.250 17.050 9.050 ;
        RECT 26.800 7.500 27.400 9.050 ;
        RECT 16.450 8.450 27.400 9.050 ;
        RECT 25.450 5.950 32.050 6.550 ;
        RECT 25.450 5.950 26.050 7.750 ;
        RECT 12.050 7.150 26.050 7.750 ;
        RECT 12.050 7.150 12.650 8.100 ;
  END 
END sdffps_6

MACRO sdffps_4
  CLASS  CORE ;
  FOREIGN sdffps_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 27.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN sb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 8.350 1.750 9.150 ;
    END
  END sb
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 21.550 9.700 23.550 10.300 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 2.700 0.000 3.300 2.700 ;
        RECT 0.000 0.000 27.500 2.500 ;
        RECT 23.750 0.000 24.350 2.700 ;
        RECT 20.600 0.000 21.200 3.750 ;
        RECT 17.950 0.000 18.550 2.650 ;
        RECT 16.850 0.000 17.450 2.650 ;
        RECT 15.750 0.000 16.350 2.650 ;
        RECT 11.550 0.000 12.150 2.800 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.100 5.950 4.100 6.550 ;
    END
  END d
  PIN se
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.350 3.450 4.350 4.050 ;
    END
  END se
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 27.500 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 18.900 9.700 20.900 10.300 ;
    END
  END qb
  PIN sdi
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.350 8.400 7.000 10.300 ;
        RECT 5.950 9.700 7.000 10.300 ;
    END
  END sdi
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 26.650 6.950 27.250 10.300 ;
        RECT 25.950 9.700 27.250 10.300 ;
    END
  END ck
  OBS 
      LAYER Metal1 ;
        RECT 1.000 5.950 1.600 7.850 ;
        RECT 1.000 7.250 4.550 7.850 ;
        RECT 2.700 7.250 4.550 7.900 ;
        RECT 2.700 7.250 3.300 9.600 ;
        RECT 7.350 7.000 8.150 7.900 ;
        RECT 5.050 7.300 8.150 7.900 ;
        RECT 5.050 7.300 5.650 9.000 ;
        RECT 4.400 8.400 5.650 9.000 ;
        RECT 7.550 7.000 8.150 9.950 ;
        RECT 4.400 8.400 5.000 9.600 ;
        RECT 7.550 9.350 8.400 9.950 ;
        RECT 8.650 5.850 11.600 6.450 ;
        RECT 8.650 5.850 9.250 8.850 ;
        RECT 8.900 8.250 9.500 9.900 ;
        RECT 8.900 9.300 10.350 9.900 ;
        RECT 16.450 6.950 21.350 7.550 ;
        RECT 16.450 6.950 17.050 8.050 ;
        RECT 12.100 5.850 24.900 6.450 ;
        RECT 12.100 5.850 12.700 7.700 ;
        RECT 9.750 7.100 12.700 7.700 ;
        RECT 24.300 5.850 24.900 7.950 ;
        RECT 14.900 5.850 15.500 8.700 ;
        RECT 25.400 5.850 26.050 6.450 ;
        RECT 10.000 8.200 14.300 8.800 ;
        RECT 11.550 8.200 14.300 8.850 ;
        RECT 25.400 5.850 26.000 9.050 ;
        RECT 17.550 8.450 26.000 9.050 ;
        RECT 13.700 7.850 14.300 10.400 ;
        RECT 17.550 8.450 18.150 10.400 ;
        RECT 13.700 9.800 18.150 10.400 ;
  END 
END sdffps_4

MACRO sdffps_3
  CLASS  CORE ;
  FOREIGN sdffps_3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 27.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN sb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 8.350 1.750 9.150 ;
    END
  END sb
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 22.150 4.700 22.800 6.200 ;
        RECT 21.800 4.700 23.300 5.300 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 27.500 2.500 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.200 5.950 4.200 6.550 ;
    END
  END d
  PIN se
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.500 4.700 5.550 5.300 ;
    END
  END se
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 27.500 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 16.850 4.700 18.850 5.300 ;
    END
  END qb
  PIN sdi
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.650 8.400 7.350 10.300 ;
        RECT 5.850 9.700 7.350 10.300 ;
    END
  END sdi
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 25.900 4.700 27.250 5.300 ;
        RECT 26.650 4.700 27.250 8.300 ;
    END
  END ck
  OBS 
      LAYER Metal1 ;
        RECT 1.000 6.650 1.600 7.850 ;
        RECT 1.000 7.250 5.000 7.850 ;
        RECT 2.700 7.250 5.000 7.900 ;
        RECT 2.700 7.250 3.300 10.350 ;
        RECT 5.550 7.300 8.450 7.900 ;
        RECT 5.550 7.300 6.150 9.000 ;
        RECT 4.400 8.400 6.150 9.000 ;
        RECT 4.400 8.400 5.000 9.600 ;
        RECT 7.850 6.300 8.450 10.300 ;
        RECT 8.950 5.850 10.400 6.450 ;
        RECT 8.950 5.850 9.550 10.350 ;
        RECT 8.950 9.750 10.700 10.350 ;
        RECT 15.350 5.300 15.950 6.500 ;
        RECT 15.350 5.900 16.700 6.500 ;
        RECT 16.100 5.900 16.700 7.600 ;
        RECT 16.100 7.000 20.250 7.600 ;
        RECT 19.650 7.600 21.500 8.200 ;
        RECT 10.750 7.150 15.600 7.750 ;
        RECT 10.750 7.150 11.350 8.050 ;
        RECT 15.000 7.150 15.600 9.300 ;
        RECT 17.300 8.100 17.900 9.300 ;
        RECT 24.150 7.350 24.750 9.300 ;
        RECT 15.000 8.700 24.750 9.300 ;
        RECT 25.550 6.350 26.150 9.450 ;
        RECT 12.050 8.250 14.500 9.150 ;
        RECT 10.050 8.550 14.500 9.150 ;
        RECT 25.500 8.850 26.300 9.450 ;
        RECT 13.900 8.250 14.500 10.400 ;
        RECT 25.500 8.850 26.100 10.400 ;
        RECT 13.900 9.800 26.100 10.400 ;
  END 
END sdffps_3

MACRO sdffps_2
  CLASS  CORE ;
  FOREIGN sdffps_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 26.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN sb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 8.350 1.750 9.150 ;
    END
  END sb
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 20.450 5.950 22.450 6.550 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 6.600 0.000 7.200 2.700 ;
        RECT 0.000 0.000 26.250 2.500 ;
        RECT 19.500 0.000 20.100 3.800 ;
        RECT 11.700 0.000 12.300 2.800 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.100 5.800 3.500 6.700 ;
    END
  END d
  PIN se
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.600 4.700 5.600 5.300 ;
    END
  END se
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 1.000 13.550 1.600 16.250 ;
        RECT 0.000 13.750 26.250 16.250 ;
        RECT 19.600 13.550 20.200 16.250 ;
        RECT 12.650 13.550 13.250 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 17.750 5.950 19.750 6.550 ;
    END
  END qb
  PIN sdi
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.200 8.450 8.200 9.050 ;
    END
  END sdi
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 24.000 7.200 26.000 7.800 ;
    END
  END ck
  OBS 
      LAYER Metal1 ;
        RECT 1.000 6.650 1.600 7.850 ;
        RECT 4.000 6.700 4.600 7.850 ;
        RECT 1.000 7.250 4.600 7.850 ;
        RECT 2.700 7.250 3.300 9.200 ;
        RECT 5.700 6.900 6.300 7.850 ;
        RECT 5.100 7.250 8.100 7.850 ;
        RECT 5.100 7.250 5.700 9.200 ;
        RECT 4.400 8.600 5.700 9.200 ;
        RECT 9.800 5.050 15.300 5.650 ;
        RECT 9.800 5.050 10.400 7.000 ;
        RECT 8.750 6.400 10.400 7.000 ;
        RECT 8.750 6.400 9.350 9.200 ;
        RECT 8.750 8.600 10.600 9.200 ;
        RECT 12.450 6.150 15.300 6.750 ;
        RECT 11.750 6.400 13.050 7.000 ;
        RECT 14.700 6.150 15.300 7.950 ;
        RECT 16.500 5.250 17.100 7.950 ;
        RECT 14.700 7.350 23.500 7.950 ;
        RECT 9.850 7.500 14.150 8.100 ;
        RECT 13.550 7.250 14.150 9.050 ;
        RECT 13.550 8.450 24.800 9.050 ;
  END 
END sdffps_2

MACRO sdffps_1
  CLASS  CORE ;
  FOREIGN sdffps_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 26.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN sb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 8.350 1.750 9.150 ;
    END
  END sb
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 20.250 5.950 22.250 6.550 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 6.600 0.000 7.200 2.700 ;
        RECT 0.000 0.000 26.250 2.500 ;
        RECT 22.300 0.000 22.900 2.600 ;
        RECT 19.300 0.000 19.900 3.750 ;
        RECT 11.700 0.000 12.300 2.800 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.100 5.800 3.500 6.700 ;
    END
  END d
  PIN se
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.400 4.700 5.400 5.300 ;
    END
  END se
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 1.000 13.550 1.600 16.250 ;
        RECT 0.000 13.750 26.250 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 17.600 5.950 19.600 6.550 ;
    END
  END qb
  PIN sdi
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.200 8.450 8.200 9.050 ;
    END
  END sdi
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 24.000 7.200 26.000 7.800 ;
    END
  END ck
  OBS 
      LAYER Metal1 ;
        RECT 1.000 6.650 1.600 7.850 ;
        RECT 4.000 6.700 4.600 7.850 ;
        RECT 1.000 7.250 4.600 7.850 ;
        RECT 2.700 7.250 3.300 9.200 ;
        RECT 5.700 6.900 6.300 7.850 ;
        RECT 5.100 7.250 8.100 7.850 ;
        RECT 5.100 7.250 5.700 9.200 ;
        RECT 4.400 8.600 5.700 9.200 ;
        RECT 9.800 5.050 15.300 5.650 ;
        RECT 9.800 5.050 10.400 7.000 ;
        RECT 8.750 6.400 10.400 7.000 ;
        RECT 8.750 6.400 9.350 9.200 ;
        RECT 8.750 8.600 10.600 9.200 ;
        RECT 12.450 6.150 15.250 6.750 ;
        RECT 11.750 6.400 13.050 7.000 ;
        RECT 14.650 6.150 15.250 7.950 ;
        RECT 16.500 5.250 17.100 7.950 ;
        RECT 14.650 7.350 23.500 7.950 ;
        RECT 9.850 7.500 14.150 8.100 ;
        RECT 13.550 7.250 14.150 9.050 ;
        RECT 13.550 8.450 24.800 9.050 ;
  END 
END sdffps_1

MACRO sdffprs_8
  CLASS  CORE ;
  FOREIGN sdffprs_8 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 37.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN sb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 25.950 8.450 26.550 10.350 ;
        RECT 17.250 9.750 26.550 10.350 ;
    END
  END sb
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 30.900 9.700 32.900 10.300 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 16.850 0.000 17.450 2.800 ;
        RECT 0.000 0.000 37.500 2.500 ;
        RECT 26.750 0.000 27.350 2.800 ;
        RECT 18.650 0.000 19.250 2.800 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.100 8.400 6.000 9.100 ;
    END
  END d
  PIN se
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.400 7.050 6.350 7.800 ;
        RECT 1.800 7.200 6.350 7.800 ;
    END
  END se
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 5.800 13.450 6.400 16.250 ;
        RECT 0.000 13.750 37.500 16.250 ;
        RECT 16.850 13.450 17.450 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 28.000 9.700 30.000 10.300 ;
    END
  END qb
  PIN sdi
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 9.400 1.650 10.300 ;
    END
  END sdi
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 35.100 7.200 37.150 7.800 ;
    END
  END ck
  PIN rb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.900 4.550 5.950 5.300 ;
        RECT 16.050 5.950 16.650 6.900 ;
        RECT 9.700 5.950 16.650 6.550 ;
        RECT 10.300 9.700 12.000 10.300 ;
        RECT 10.300 8.550 10.900 10.300 ;
        RECT 9.700 4.700 10.300 9.150 ;
        RECT 4.900 4.700 10.300 5.300 ;
    END
  END rb
  OBS 
      LAYER Metal1 ;
        RECT 1.950 5.950 7.850 6.550 ;
        RECT 2.150 9.700 9.750 10.300 ;
        RECT 18.550 7.550 20.850 8.150 ;
        RECT 12.850 4.700 25.550 5.300 ;
        RECT 24.950 4.800 31.150 5.400 ;
        RECT 33.950 5.850 34.550 7.800 ;
        RECT 23.450 7.200 34.550 7.800 ;
        RECT 11.850 8.500 14.850 9.100 ;
        RECT 23.450 7.200 24.050 9.250 ;
        RECT 14.250 8.650 24.050 9.250 ;
        RECT 14.250 8.500 14.850 10.200 ;
        RECT 32.250 4.700 35.850 5.300 ;
        RECT 32.250 4.700 32.850 6.600 ;
        RECT 17.150 6.000 32.850 6.600 ;
        RECT 17.150 6.000 17.750 8.000 ;
        RECT 11.050 7.400 17.750 8.000 ;
        RECT 22.050 6.000 22.650 8.150 ;
  END 
END sdffprs_8

MACRO sdffprs_6
  CLASS  CORE ;
  FOREIGN sdffprs_6 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 36.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN sb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 24.700 8.450 25.300 10.300 ;
        RECT 24.700 8.450 26.550 9.050 ;
        RECT 17.100 9.700 25.300 10.300 ;
    END
  END sb
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 30.050 9.700 32.050 10.300 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 16.800 0.000 17.400 2.800 ;
        RECT 0.000 0.000 36.250 2.500 ;
        RECT 25.800 0.000 26.400 2.800 ;
        RECT 18.500 0.000 19.100 2.800 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.150 8.450 6.150 9.050 ;
    END
  END d
  PIN se
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.200 7.200 6.550 7.800 ;
    END
  END se
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 6.000 13.450 6.600 16.250 ;
        RECT 0.000 13.750 36.250 16.250 ;
        RECT 16.700 13.450 17.300 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 27.350 9.700 29.350 10.300 ;
    END
  END qb
  PIN sdi
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 9.550 1.750 10.450 ;
    END
  END sdi
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 33.900 7.200 35.900 7.800 ;
    END
  END ck
  PIN rb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.450 4.700 10.300 5.300 ;
        RECT 16.050 5.950 16.650 6.900 ;
        RECT 9.550 5.950 16.650 6.550 ;
        RECT 10.050 9.800 11.350 10.400 ;
        RECT 10.050 8.600 10.650 10.400 ;
        RECT 9.550 4.700 10.300 6.550 ;
        RECT 9.550 4.700 10.150 9.200 ;
        RECT 9.150 4.700 10.300 5.400 ;
    END
  END rb
  OBS 
      LAYER Metal1 ;
        RECT 2.350 5.950 7.850 6.550 ;
        RECT 2.250 9.700 9.550 10.300 ;
        RECT 18.700 7.450 21.000 8.050 ;
        RECT 18.700 7.450 19.300 8.100 ;
        RECT 12.900 4.700 30.200 5.300 ;
        RECT 24.050 4.700 24.650 5.450 ;
        RECT 23.300 7.200 33.350 7.800 ;
        RECT 23.300 7.200 23.900 9.200 ;
        RECT 11.650 8.600 23.900 9.200 ;
        RECT 14.250 8.600 14.850 9.250 ;
        RECT 11.650 8.600 12.250 9.300 ;
        RECT 17.200 5.950 34.600 6.550 ;
        RECT 10.650 7.200 15.550 7.800 ;
        RECT 22.200 5.950 22.800 7.850 ;
        RECT 17.200 5.950 17.800 8.050 ;
        RECT 14.950 7.400 17.800 8.050 ;
  END 
END sdffprs_6

MACRO sdffprs_4
  CLASS  CORE ;
  FOREIGN sdffprs_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 32.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN sb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 18.900 9.350 19.700 10.300 ;
        RECT 18.900 9.600 20.800 10.300 ;
    END
  END sb
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 26.050 9.700 28.050 10.300 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 15.200 0.000 15.900 2.800 ;
        RECT 0.000 0.000 32.500 2.500 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 8.350 1.750 9.150 ;
    END
  END d
  PIN se
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.450 5.900 3.250 6.600 ;
    END
  END se
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.450 13.500 1.050 16.250 ;
        RECT 0.000 13.750 32.500 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 22.550 9.700 24.550 10.300 ;
    END
  END qb
  PIN sdi
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.250 9.700 7.250 10.300 ;
    END
  END sdi
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 30.950 4.700 32.250 5.300 ;
        RECT 31.650 4.700 32.250 8.200 ;
    END
  END ck
  PIN rb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.050 4.700 7.800 5.300 ;
        RECT 14.450 5.950 15.050 7.000 ;
        RECT 7.200 5.950 15.050 6.550 ;
        RECT 7.200 4.700 7.800 6.550 ;
    END
  END rb
  OBS 
      LAYER Metal1 ;
        RECT 0.350 6.850 0.950 7.850 ;
        RECT 3.750 6.900 4.350 7.850 ;
        RECT 0.350 7.250 4.350 7.850 ;
        RECT 2.250 7.250 2.850 9.200 ;
        RECT 5.450 6.750 6.050 7.850 ;
        RECT 4.850 7.250 7.750 7.850 ;
        RECT 4.850 7.250 5.450 9.050 ;
        RECT 3.950 8.450 5.450 9.050 ;
        RECT 15.550 9.800 18.400 10.400 ;
        RECT 11.000 4.850 26.600 5.450 ;
        RECT 26.000 4.850 26.600 6.850 ;
        RECT 16.150 6.000 24.950 6.600 ;
        RECT 21.150 6.000 21.750 6.900 ;
        RECT 24.200 6.000 24.950 7.950 ;
        RECT 8.450 7.300 13.350 7.900 ;
        RECT 8.450 7.300 9.050 7.950 ;
        RECT 29.100 6.450 29.700 7.950 ;
        RECT 24.200 7.350 29.700 7.950 ;
        RECT 16.150 6.000 16.750 8.200 ;
        RECT 12.750 7.600 16.750 8.200 ;
        RECT 12.750 7.300 13.350 9.300 ;
        RECT 30.400 5.900 31.050 6.500 ;
        RECT 22.800 7.500 23.400 9.050 ;
        RECT 17.650 8.250 23.400 8.850 ;
        RECT 21.150 8.450 31.000 9.050 ;
        RECT 14.400 8.700 18.250 9.300 ;
        RECT 30.400 5.900 31.000 9.950 ;
        RECT 30.400 9.350 31.300 9.950 ;
        RECT 14.400 8.700 15.000 10.400 ;
        RECT 8.450 9.800 15.000 10.400 ;
  END 
END sdffprs_4

MACRO sdffprs_3
  CLASS  CORE ;
  FOREIGN sdffprs_3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 31.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN sb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 18.900 9.350 19.700 10.300 ;
        RECT 18.900 9.600 20.800 10.300 ;
    END
  END sb
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 25.050 9.700 27.050 10.300 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 15.250 0.000 15.850 2.800 ;
        RECT 0.000 0.000 31.250 2.500 ;
        RECT 17.250 0.000 17.850 2.700 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 8.350 1.750 9.150 ;
    END
  END d
  PIN se
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.450 5.900 3.250 6.600 ;
    END
  END se
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.450 13.500 1.050 16.250 ;
        RECT 0.000 13.750 31.250 16.250 ;
        RECT 20.950 13.550 21.550 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 22.050 9.700 24.050 10.300 ;
    END
  END qb
  PIN sdi
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.250 9.700 7.250 10.300 ;
    END
  END sdi
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 29.700 4.700 31.000 5.300 ;
        RECT 30.400 4.700 31.000 8.200 ;
    END
  END ck
  PIN rb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.050 4.700 7.800 5.300 ;
        RECT 14.150 5.950 14.750 6.800 ;
        RECT 7.200 5.950 14.750 6.550 ;
        RECT 7.200 4.700 7.800 6.550 ;
    END
  END rb
  OBS 
      LAYER Metal1 ;
        RECT 0.350 6.850 0.950 7.850 ;
        RECT 3.750 6.900 4.350 7.850 ;
        RECT 0.350 7.250 4.350 7.850 ;
        RECT 2.250 7.250 2.850 9.200 ;
        RECT 5.450 6.700 6.050 7.850 ;
        RECT 4.850 7.250 7.750 7.850 ;
        RECT 4.850 7.250 5.450 9.050 ;
        RECT 3.950 8.450 5.450 9.050 ;
        RECT 15.350 9.600 18.400 10.300 ;
        RECT 11.050 4.600 20.950 5.200 ;
        RECT 11.050 4.600 11.650 5.450 ;
        RECT 20.250 6.950 25.350 7.550 ;
        RECT 24.750 6.950 25.350 7.950 ;
        RECT 16.500 5.850 28.500 6.450 ;
        RECT 16.500 5.850 17.100 7.900 ;
        RECT 8.250 7.300 17.100 7.900 ;
        RECT 27.900 5.850 28.500 7.950 ;
        RECT 13.150 7.300 13.750 9.300 ;
        RECT 17.800 8.050 22.150 8.850 ;
        RECT 14.250 8.400 18.400 9.000 ;
        RECT 8.250 8.450 12.200 9.050 ;
        RECT 21.550 8.450 29.900 9.050 ;
        RECT 29.300 6.250 29.900 10.050 ;
        RECT 11.600 8.450 12.200 10.400 ;
        RECT 29.300 9.450 30.250 10.050 ;
        RECT 14.250 8.400 14.850 10.400 ;
        RECT 11.600 9.800 14.850 10.400 ;
  END 
END sdffprs_3

MACRO sdffprs_2
  CLASS  CORE ;
  FOREIGN sdffprs_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 31.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN sb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 18.450 9.700 20.450 10.300 ;
    END
  END sb
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 25.250 9.700 27.250 10.300 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 15.100 0.000 15.700 2.700 ;
        RECT 0.000 0.000 31.250 2.500 ;
        RECT 17.550 0.000 18.150 2.700 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.350 8.350 1.850 9.150 ;
    END
  END d
  PIN se
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.250 5.950 3.250 6.550 ;
    END
  END se
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.500 13.600 1.100 16.250 ;
        RECT 0.000 13.750 31.250 16.250 ;
        RECT 19.050 13.550 19.650 16.250 ;
        RECT 15.600 13.550 16.200 16.250 ;
        RECT 4.600 13.550 5.200 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 21.850 9.700 23.850 10.300 ;
    END
  END qb
  PIN sdi
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.250 9.700 7.250 10.300 ;
    END
  END sdi
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 30.300 6.650 30.900 7.800 ;
        RECT 29.000 7.200 31.000 7.800 ;
    END
  END ck
  PIN rb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.050 4.700 7.800 5.300 ;
        RECT 7.200 5.950 10.400 6.550 ;
        RECT 7.200 4.700 7.800 6.550 ;
    END
  END rb
  OBS 
      LAYER Metal1 ;
        RECT 3.750 6.900 4.350 7.850 ;
        RECT 0.350 7.250 4.350 7.850 ;
        RECT 2.350 7.250 2.950 9.200 ;
        RECT 5.450 6.700 6.050 7.850 ;
        RECT 4.850 7.250 7.800 7.850 ;
        RECT 4.850 7.250 5.450 9.050 ;
        RECT 4.050 8.450 5.450 9.050 ;
        RECT 10.400 3.450 16.850 4.050 ;
        RECT 15.100 9.750 17.950 10.350 ;
        RECT 16.250 7.350 25.250 7.950 ;
        RECT 12.650 7.550 16.850 8.150 ;
        RECT 12.650 7.550 13.250 8.850 ;
        RECT 10.900 8.250 13.250 8.850 ;
        RECT 15.150 6.250 28.300 6.850 ;
        RECT 10.900 6.450 15.750 7.050 ;
        RECT 10.900 6.450 11.500 7.750 ;
        RECT 8.500 7.150 11.500 7.750 ;
        RECT 27.700 6.250 28.300 7.800 ;
        RECT 17.350 8.450 29.950 9.050 ;
        RECT 14.000 8.650 17.950 9.250 ;
        RECT 14.000 8.650 14.600 9.950 ;
        RECT 8.500 9.350 14.600 9.950 ;
  END 
END sdffprs_2

MACRO sdffprs_1
  CLASS  CORE ;
  FOREIGN sdffprs_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 31.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN sb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 18.450 9.650 20.400 10.300 ;
    END
  END sb
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 25.050 9.700 27.050 10.300 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 15.100 0.000 15.700 2.700 ;
        RECT 0.000 0.000 31.250 2.500 ;
        RECT 17.550 0.000 18.150 2.700 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.350 8.350 1.850 9.150 ;
    END
  END d
  PIN se
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.250 5.950 3.250 6.550 ;
    END
  END se
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.500 13.600 1.100 16.250 ;
        RECT 0.000 13.750 31.250 16.250 ;
        RECT 19.050 13.550 19.650 16.250 ;
        RECT 15.600 13.550 16.200 16.250 ;
        RECT 4.600 13.550 5.200 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 21.850 9.700 23.850 10.300 ;
    END
  END qb
  PIN sdi
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.250 9.700 7.250 10.300 ;
    END
  END sdi
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 29.000 7.200 31.000 7.800 ;
    END
  END ck
  PIN rb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.050 4.700 7.800 5.300 ;
        RECT 7.200 5.950 10.400 6.550 ;
        RECT 7.200 4.700 7.800 6.550 ;
    END
  END rb
  OBS 
      LAYER Metal1 ;
        RECT 3.750 6.900 4.350 7.850 ;
        RECT 0.350 7.250 4.350 7.850 ;
        RECT 2.350 7.250 2.950 9.200 ;
        RECT 5.450 6.750 6.050 7.850 ;
        RECT 4.850 7.250 7.800 7.850 ;
        RECT 4.850 7.250 5.450 9.050 ;
        RECT 4.050 8.450 5.450 9.050 ;
        RECT 10.400 3.450 16.850 4.050 ;
        RECT 15.100 9.750 17.950 10.350 ;
        RECT 16.250 7.350 25.250 7.950 ;
        RECT 12.650 7.550 16.850 8.150 ;
        RECT 12.650 7.550 13.250 8.850 ;
        RECT 10.900 8.250 13.250 8.850 ;
        RECT 15.150 6.250 28.300 6.850 ;
        RECT 10.900 6.450 15.750 7.050 ;
        RECT 10.900 6.450 11.500 7.750 ;
        RECT 8.500 7.150 11.500 7.750 ;
        RECT 27.700 6.250 28.300 7.800 ;
        RECT 17.350 8.450 29.600 9.050 ;
        RECT 14.000 8.650 17.950 9.250 ;
        RECT 14.000 8.650 14.600 9.950 ;
        RECT 8.500 9.350 14.600 9.950 ;
  END 
END sdffprs_1

MACRO sdffpr_8
  CLASS  CORE ;
  FOREIGN sdffpr_8 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 35.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 23.600 9.700 27.600 10.300 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 22.300 0.000 22.900 2.800 ;
        RECT 0.000 0.000 35.000 2.500 ;
        RECT 32.100 0.000 32.700 2.800 ;
        RECT 25.300 0.000 25.900 2.800 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.550 4.700 5.150 5.300 ;
    END
  END d
  PIN se
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.650 8.350 7.700 9.050 ;
        RECT 1.600 8.450 7.700 9.050 ;
        RECT 7.100 7.900 7.700 9.050 ;
    END
  END se
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 1.000 13.450 1.600 16.250 ;
        RECT 0.000 13.750 35.000 16.250 ;
        RECT 32.100 13.450 32.700 16.250 ;
        RECT 25.300 13.450 25.900 16.250 ;
        RECT 20.600 13.450 21.200 16.250 ;
        RECT 4.800 13.450 5.400 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 29.550 8.450 31.550 9.050 ;
    END
  END qb
  PIN sdi
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.350 4.700 8.350 5.300 ;
    END
  END sdi
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 32.500 4.700 34.500 5.300 ;
    END
  END ck
  PIN rb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.350 4.700 2.050 5.450 ;
    END
  END rb
  OBS 
      LAYER Metal1 ;
        RECT 1.600 7.150 6.400 7.750 ;
        RECT 1.450 5.950 8.800 6.550 ;
        RECT 8.200 6.200 9.550 6.800 ;
        RECT 8.200 5.950 8.800 10.300 ;
        RECT 1.000 9.700 8.800 10.300 ;
        RECT 10.050 5.100 11.250 5.700 ;
        RECT 10.050 5.100 10.650 10.300 ;
        RECT 10.050 9.700 10.700 10.300 ;
        RECT 15.150 6.100 19.150 6.700 ;
        RECT 11.650 6.250 15.750 6.850 ;
        RECT 11.650 6.250 12.250 9.050 ;
        RECT 11.150 8.450 16.550 9.050 ;
        RECT 14.050 5.000 21.100 5.600 ;
        RECT 14.050 5.000 14.650 5.750 ;
        RECT 20.500 5.000 21.100 6.650 ;
        RECT 14.650 9.550 15.250 10.250 ;
        RECT 14.650 9.650 22.900 10.250 ;
        RECT 22.500 8.450 26.250 9.050 ;
        RECT 17.250 8.550 23.100 9.150 ;
        RECT 24.000 5.300 29.700 5.900 ;
        RECT 21.400 7.200 34.400 7.800 ;
        RECT 12.750 7.350 22.000 7.950 ;
  END 
END sdffpr_8

MACRO sdffpr_6
  CLASS  CORE ;
  FOREIGN sdffpr_6 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 33.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 28.250 9.700 30.350 10.300 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 16.700 0.000 17.300 2.800 ;
        RECT 0.000 0.000 33.750 2.500 ;
        RECT 30.950 0.000 31.550 2.800 ;
        RECT 27.550 0.000 28.150 2.800 ;
        RECT 22.850 0.000 23.450 2.800 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.450 4.700 5.250 5.400 ;
    END
  END d
  PIN se
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.250 7.650 7.850 9.050 ;
        RECT 2.100 8.450 7.850 9.050 ;
    END
  END se
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 1.250 13.450 1.850 16.250 ;
        RECT 0.000 13.750 33.750 16.250 ;
        RECT 27.550 13.450 28.150 16.250 ;
        RECT 24.550 13.450 25.150 16.250 ;
        RECT 21.150 13.450 21.750 16.250 ;
        RECT 5.450 13.450 6.050 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 22.350 5.950 25.150 6.550 ;
    END
  END qb
  PIN sdi
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.550 4.700 8.600 5.300 ;
    END
  END sdi
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 31.250 4.700 33.250 5.300 ;
    END
  END ck
  PIN rb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.400 4.700 2.200 5.400 ;
    END
  END rb
  OBS 
      LAYER Metal1 ;
        RECT 2.250 7.150 6.550 7.750 ;
        RECT 1.000 5.900 9.650 6.500 ;
        RECT 8.550 5.900 9.150 10.300 ;
        RECT 1.100 9.700 9.150 10.300 ;
        RECT 10.150 5.150 11.350 5.750 ;
        RECT 10.150 5.150 10.750 7.900 ;
        RECT 9.650 7.300 10.250 10.350 ;
        RECT 9.650 9.750 10.950 10.350 ;
        RECT 11.250 6.250 19.950 6.850 ;
        RECT 11.250 6.250 11.850 9.250 ;
        RECT 13.550 8.450 17.200 9.050 ;
        RECT 10.750 8.650 14.150 9.250 ;
        RECT 14.350 5.150 21.600 5.750 ;
        RECT 21.000 5.150 21.600 6.850 ;
        RECT 15.300 9.650 26.450 10.250 ;
        RECT 17.900 8.450 31.150 9.050 ;
        RECT 12.350 7.350 33.300 7.950 ;
        RECT 12.350 7.350 12.950 8.150 ;
  END 
END sdffpr_6

MACRO sdffpr_4
  CLASS  CORE ;
  FOREIGN sdffpr_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 28.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 22.300 5.950 24.300 6.550 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 28.750 2.500 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.100 4.700 2.800 5.450 ;
    END
  END d
  PIN se
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.500 4.700 5.500 5.300 ;
    END
  END se
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 28.750 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 19.300 5.950 21.300 6.550 ;
    END
  END qb
  PIN sdi
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.650 8.400 7.300 10.300 ;
        RECT 5.850 9.700 7.300 10.300 ;
    END
  END sdi
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 27.200 4.700 28.500 5.300 ;
        RECT 27.900 4.700 28.500 7.650 ;
    END
  END ck
  PIN rb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.950 7.200 1.550 9.050 ;
        RECT 0.950 7.200 2.900 7.800 ;
        RECT 0.350 8.450 1.550 9.050 ;
    END
  END rb
  OBS 
      LAYER Metal1 ;
        RECT 0.300 5.950 4.050 6.550 ;
        RECT 3.450 7.300 5.000 7.900 ;
        RECT 3.450 5.950 4.050 9.250 ;
        RECT 2.700 8.650 4.050 9.250 ;
        RECT 5.550 7.300 9.150 7.900 ;
        RECT 5.550 7.300 6.150 9.000 ;
        RECT 4.600 8.400 6.150 9.000 ;
        RECT 4.600 8.400 5.200 9.600 ;
        RECT 16.350 5.850 16.950 6.500 ;
        RECT 9.650 5.900 16.950 6.500 ;
        RECT 9.650 5.900 10.250 10.300 ;
        RECT 9.650 9.700 11.350 10.300 ;
        RECT 10.800 7.200 11.400 7.950 ;
        RECT 25.550 6.450 26.150 7.950 ;
        RECT 10.800 7.350 26.150 7.950 ;
        RECT 15.600 7.350 16.200 9.050 ;
        RECT 26.800 5.900 27.400 9.700 ;
        RECT 20.050 8.450 27.400 9.050 ;
        RECT 10.750 8.600 14.300 9.200 ;
        RECT 26.800 9.000 27.550 9.700 ;
        RECT 13.700 8.450 14.300 10.400 ;
        RECT 18.550 9.300 20.650 9.900 ;
        RECT 20.050 8.450 20.650 9.900 ;
        RECT 13.700 9.800 19.150 10.400 ;
  END 
END sdffpr_4

MACRO sdffpr_3
  CLASS  CORE ;
  FOREIGN sdffpr_3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 27.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 21.300 5.950 23.300 6.550 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 27.500 2.500 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.150 4.700 1.750 6.000 ;
        RECT 1.150 4.700 2.900 5.400 ;
    END
  END d
  PIN se
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.350 8.100 3.950 9.100 ;
        RECT 4.000 9.700 5.400 10.300 ;
        RECT 4.000 8.500 4.600 10.300 ;
        RECT 3.350 8.500 4.600 9.100 ;
    END
  END se
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 27.500 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 18.750 5.950 20.750 6.550 ;
    END
  END qb
  PIN sdi
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.700 8.400 7.300 10.300 ;
        RECT 6.700 9.700 7.950 10.300 ;
    END
  END sdi
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 25.950 4.700 27.250 5.300 ;
        RECT 26.650 4.700 27.250 8.350 ;
    END
  END ck
  PIN rb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.450 7.550 1.050 9.050 ;
        RECT 0.450 8.450 1.700 9.050 ;
    END
  END rb
  OBS 
      LAYER Metal1 ;
        RECT 2.450 5.900 6.850 6.550 ;
        RECT 2.450 5.900 3.050 7.400 ;
        RECT 2.200 6.800 2.800 10.400 ;
        RECT 2.200 9.800 3.300 10.400 ;
        RECT 4.550 7.200 8.550 7.800 ;
        RECT 9.050 4.900 16.350 5.500 ;
        RECT 15.750 4.900 16.350 5.600 ;
        RECT 9.050 4.900 9.650 10.450 ;
        RECT 9.050 9.850 10.950 10.450 ;
        RECT 10.700 6.350 18.050 6.950 ;
        RECT 17.450 6.350 18.050 7.950 ;
        RECT 10.700 6.350 11.300 7.900 ;
        RECT 17.450 7.350 24.750 7.950 ;
        RECT 15.350 6.350 15.950 9.200 ;
        RECT 10.150 8.450 10.750 9.200 ;
        RECT 17.600 8.450 26.150 9.050 ;
        RECT 13.400 7.500 14.050 9.200 ;
        RECT 10.150 8.600 14.050 9.200 ;
        RECT 25.550 6.450 26.150 9.900 ;
        RECT 13.400 7.500 14.000 10.350 ;
        RECT 25.550 9.300 26.300 9.900 ;
        RECT 17.600 8.450 18.200 10.350 ;
        RECT 13.400 9.750 18.200 10.350 ;
  END 
END sdffpr_3

MACRO sdffpr_2
  CLASS  CORE ;
  FOREIGN sdffpr_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 26.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 20.750 5.950 22.750 6.550 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 11.300 0.000 11.900 2.700 ;
        RECT 0.000 0.000 26.250 2.500 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.100 5.950 4.100 6.550 ;
    END
  END d
  PIN se
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.500 3.450 4.500 4.050 ;
    END
  END se
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 1.000 13.550 1.600 16.250 ;
        RECT 0.000 13.750 26.250 16.250 ;
        RECT 19.450 13.450 20.050 16.250 ;
        RECT 9.350 13.450 9.950 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 17.900 5.950 19.900 6.550 ;
    END
  END qb
  PIN sdi
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.400 8.350 7.900 9.150 ;
    END
  END sdi
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 24.000 8.450 26.000 9.050 ;
    END
  END ck
  PIN rb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 8.350 1.750 9.150 ;
    END
  END rb
  OBS 
      LAYER Metal1 ;
        RECT 1.000 6.900 1.600 7.850 ;
        RECT 1.000 7.250 4.700 7.850 ;
        RECT 2.400 7.250 3.000 9.200 ;
        RECT 6.550 5.300 8.100 5.900 ;
        RECT 6.550 5.300 7.150 6.950 ;
        RECT 5.200 6.350 7.150 6.950 ;
        RECT 5.200 6.350 5.800 9.050 ;
        RECT 4.100 8.450 5.800 9.050 ;
        RECT 8.900 5.800 15.400 6.400 ;
        RECT 8.400 6.400 9.500 7.000 ;
        RECT 8.400 6.400 9.000 9.200 ;
        RECT 8.400 8.600 10.500 9.200 ;
        RECT 11.100 8.450 23.500 9.050 ;
        RECT 14.300 8.450 15.000 9.200 ;
        RECT 10.000 7.200 24.800 7.800 ;
        RECT 9.500 7.500 10.600 8.100 ;
        RECT 24.450 3.200 25.050 3.950 ;
        RECT 16.600 3.350 25.050 3.950 ;
  END 
END sdffpr_2

MACRO sdffpr_1
  CLASS  CORE ;
  FOREIGN sdffpr_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 26.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 20.250 5.950 22.250 6.550 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 11.300 0.000 11.900 2.700 ;
        RECT 0.000 0.000 26.250 2.500 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.100 5.950 4.100 6.550 ;
    END
  END d
  PIN se
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.500 3.450 4.500 4.050 ;
    END
  END se
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 1.000 13.550 1.600 16.250 ;
        RECT 0.000 13.750 26.250 16.250 ;
        RECT 9.350 13.450 9.950 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 17.400 5.950 19.400 6.550 ;
    END
  END qb
  PIN sdi
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.300 8.350 7.900 9.100 ;
    END
  END sdi
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 24.000 8.450 26.000 9.050 ;
    END
  END ck
  PIN rb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 8.350 1.750 9.150 ;
    END
  END rb
  OBS 
      LAYER Metal1 ;
        RECT 1.000 6.900 1.600 7.800 ;
        RECT 1.000 7.200 4.700 7.800 ;
        RECT 2.400 7.200 3.000 9.200 ;
        RECT 6.550 5.300 8.100 5.900 ;
        RECT 6.550 5.300 7.150 6.550 ;
        RECT 5.200 5.950 7.150 6.550 ;
        RECT 5.200 5.950 5.800 9.050 ;
        RECT 4.100 8.450 5.800 9.050 ;
        RECT 8.900 5.800 15.400 6.400 ;
        RECT 8.400 6.400 9.500 7.000 ;
        RECT 8.400 6.400 9.000 9.200 ;
        RECT 8.400 8.600 10.600 9.200 ;
        RECT 11.100 8.450 23.500 9.050 ;
        RECT 14.300 8.450 15.000 9.200 ;
        RECT 10.050 7.200 24.850 7.800 ;
        RECT 9.500 7.500 10.650 8.100 ;
        RECT 24.450 3.200 25.050 3.950 ;
        RECT 16.600 3.350 25.050 3.950 ;
  END 
END sdffpr_1

MACRO sdffphc_8
  CLASS  CORE ;
  FOREIGN sdffphc_8 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 40.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 34.600 9.700 36.600 10.300 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 19.300 0.000 19.900 2.800 ;
        RECT 0.000 0.000 40.000 2.500 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.900 8.450 3.900 9.050 ;
    END
  END d
  PIN se
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.700 7.200 12.450 7.800 ;
    END
  END se
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 5.250 13.450 5.850 16.250 ;
        RECT 0.000 13.750 40.000 16.250 ;
        RECT 30.250 13.450 30.850 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 31.050 9.700 33.050 10.300 ;
    END
  END qb
  PIN g
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.300 7.100 7.050 7.800 ;
    END
  END g
  PIN sdi
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 11.000 8.450 13.000 9.050 ;
    END
  END sdi
  PIN clb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 4.700 2.250 5.300 ;
    END
  END clb
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 37.450 4.700 39.450 5.300 ;
    END
  END ck
  OBS 
      LAYER Metal1 ;
        RECT 2.150 5.950 8.900 6.550 ;
        RECT 10.050 5.950 14.250 6.550 ;
        RECT 13.650 5.950 14.250 10.450 ;
        RECT 10.050 9.850 14.250 10.450 ;
        RECT 15.350 6.100 15.950 10.350 ;
        RECT 23.650 5.900 26.000 6.500 ;
        RECT 25.400 5.700 26.000 6.500 ;
        RECT 17.600 5.950 24.250 6.550 ;
        RECT 17.600 5.950 18.200 9.050 ;
        RECT 17.600 8.450 22.950 9.050 ;
        RECT 7.750 4.550 17.100 5.150 ;
        RECT 16.500 4.550 17.100 10.300 ;
        RECT 16.500 9.700 29.150 10.300 ;
        RECT 23.450 4.600 27.550 5.200 ;
        RECT 23.450 4.600 24.050 5.250 ;
        RECT 26.950 4.650 34.650 5.250 ;
        RECT 25.400 7.000 26.000 7.800 ;
        RECT 18.900 7.200 39.350 7.800 ;
  END 
END sdffphc_8

MACRO sdffphc_6
  CLASS  CORE ;
  FOREIGN sdffphc_6 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 38.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 33.400 9.700 35.400 10.300 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 26.150 0.000 26.750 2.800 ;
        RECT 0.000 0.000 38.750 2.500 ;
        RECT 32.550 0.000 33.150 2.800 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.950 8.450 4.050 9.050 ;
    END
  END d
  PIN se
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 10.050 7.200 12.900 7.800 ;
    END
  END se
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 32.550 13.450 33.150 16.250 ;
        RECT 0.000 13.750 38.750 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 27.850 8.450 29.850 9.050 ;
    END
  END qb
  PIN g
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.700 7.050 7.350 7.800 ;
    END
  END g
  PIN sdi
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 11.750 4.700 13.750 5.300 ;
    END
  END sdi
  PIN clb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.350 5.750 1.650 6.750 ;
    END
  END clb
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 36.250 5.950 38.250 6.550 ;
    END
  END ck
  OBS 
      LAYER Metal1 ;
        RECT 2.150 5.950 9.150 6.550 ;
        RECT 10.250 5.950 14.750 6.550 ;
        RECT 14.150 5.950 14.750 10.200 ;
        RECT 10.250 9.600 14.750 10.200 ;
        RECT 15.450 4.900 16.450 5.500 ;
        RECT 15.450 4.900 16.050 10.300 ;
        RECT 15.450 9.700 16.550 10.300 ;
        RECT 16.800 5.950 24.900 6.550 ;
        RECT 16.800 5.950 17.400 9.000 ;
        RECT 16.800 8.400 21.650 9.000 ;
        RECT 19.750 9.500 20.350 10.250 ;
        RECT 19.750 9.650 31.450 10.250 ;
        RECT 26.500 7.100 32.750 7.700 ;
        RECT 26.500 7.100 27.100 9.000 ;
        RECT 22.350 8.400 27.100 9.000 ;
        RECT 25.400 6.000 34.500 6.600 ;
        RECT 33.900 6.000 34.500 7.800 ;
        RECT 33.900 7.200 38.300 7.800 ;
        RECT 25.400 6.000 26.000 7.900 ;
        RECT 17.950 7.300 26.000 7.900 ;
  END 
END sdffphc_6

MACRO sdffphc_4
  CLASS  CORE ;
  FOREIGN sdffphc_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 35.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 30.450 7.200 32.450 7.800 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 22.450 0.000 23.050 2.700 ;
        RECT 0.000 0.000 35.000 2.500 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.350 7.300 1.950 10.300 ;
        RECT 1.350 9.600 5.100 10.300 ;
        RECT 4.500 8.500 5.100 10.300 ;
    END
  END d
  PIN se
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.100 4.700 11.300 5.300 ;
    END
  END se
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 17.750 13.500 18.450 16.250 ;
        RECT 0.000 13.750 35.000 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 26.250 5.950 28.250 6.550 ;
    END
  END qb
  PIN g
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 5.950 0.850 9.600 ;
        RECT 0.250 5.950 1.550 6.550 ;
    END
  END g
  PIN sdi
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 11.800 4.700 13.800 5.300 ;
    END
  END sdi
  PIN clb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.700 4.700 8.000 5.300 ;
    END
  END clb
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 18.300 5.950 20.300 6.550 ;
    END
  END ck
  OBS 
      LAYER Metal1 ;
        RECT 2.450 5.650 5.200 6.250 ;
        RECT 4.600 5.900 7.300 6.500 ;
        RECT 6.700 5.900 7.300 7.650 ;
        RECT 9.250 6.550 9.850 7.650 ;
        RECT 6.700 7.050 9.850 7.650 ;
        RECT 2.450 5.650 3.050 9.100 ;
        RECT 2.450 8.500 4.000 9.100 ;
        RECT 8.050 7.050 8.650 9.100 ;
        RECT 10.700 6.550 11.550 7.150 ;
        RECT 10.700 6.550 11.300 9.100 ;
        RECT 10.700 8.450 13.250 9.100 ;
        RECT 9.750 8.500 13.250 9.100 ;
        RECT 14.700 5.400 16.000 6.000 ;
        RECT 14.700 5.400 15.300 7.100 ;
        RECT 13.750 6.500 15.300 7.100 ;
        RECT 13.750 6.500 14.350 9.300 ;
        RECT 13.750 8.700 15.450 9.300 ;
        RECT 14.850 7.600 16.550 8.200 ;
        RECT 15.950 7.600 16.550 9.050 ;
        RECT 15.950 8.450 25.150 9.050 ;
        RECT 15.800 6.500 17.650 7.100 ;
        RECT 17.050 6.500 17.650 7.950 ;
        RECT 17.050 7.350 25.700 7.950 ;
        RECT 3.550 6.800 4.150 7.600 ;
        RECT 3.550 7.000 6.200 7.600 ;
        RECT 5.600 7.000 6.200 10.400 ;
        RECT 28.450 8.100 29.050 10.400 ;
        RECT 5.600 9.800 29.050 10.400 ;
  END 
END sdffphc_4

MACRO sdffphc_3
  CLASS  CORE ;
  FOREIGN sdffphc_3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 32.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 28.750 5.950 30.750 6.550 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 32.500 2.500 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.450 7.350 2.050 10.300 ;
        RECT 1.450 9.550 5.100 10.300 ;
    END
  END d
  PIN se
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.950 4.700 8.550 7.100 ;
        RECT 7.950 4.700 9.050 5.300 ;
    END
  END se
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 32.500 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 25.050 5.950 27.050 6.550 ;
    END
  END qb
  PIN g
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.350 5.950 0.950 9.050 ;
        RECT 0.350 5.950 1.550 6.550 ;
    END
  END g
  PIN sdi
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 10.650 4.700 12.800 5.300 ;
    END
  END sdi
  PIN clb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.950 4.700 7.250 5.300 ;
        RECT 6.650 4.700 7.250 6.500 ;
    END
  END clb
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 18.450 5.950 20.450 6.550 ;
    END
  END ck
  OBS 
      LAYER Metal1 ;
        RECT 3.200 5.900 6.000 6.500 ;
        RECT 5.400 5.900 6.000 7.600 ;
        RECT 5.400 7.000 7.350 7.600 ;
        RECT 9.050 6.500 9.650 8.200 ;
        RECT 8.150 7.600 9.650 8.200 ;
        RECT 6.750 7.000 7.350 9.300 ;
        RECT 3.200 5.900 3.800 9.050 ;
        RECT 8.150 7.600 8.750 9.300 ;
        RECT 6.750 8.700 8.750 9.300 ;
        RECT 10.750 8.450 13.050 9.050 ;
        RECT 10.750 6.400 11.350 9.300 ;
        RECT 9.850 8.700 11.350 9.300 ;
        RECT 13.550 5.200 15.700 5.800 ;
        RECT 13.550 5.200 14.150 9.300 ;
        RECT 13.550 8.700 15.300 9.300 ;
        RECT 14.850 6.300 17.650 6.900 ;
        RECT 17.050 6.300 17.650 7.950 ;
        RECT 17.050 7.350 24.750 7.950 ;
        RECT 14.650 7.600 16.400 8.200 ;
        RECT 15.800 7.600 16.400 9.050 ;
        RECT 15.800 8.450 25.650 9.050 ;
        RECT 4.300 7.000 4.900 8.700 ;
        RECT 4.300 8.100 6.250 8.700 ;
        RECT 5.650 8.100 6.250 10.400 ;
        RECT 18.750 9.550 28.250 10.150 ;
        RECT 27.650 7.350 28.250 10.150 ;
        RECT 5.650 9.800 19.650 10.400 ;
  END 
END sdffphc_3

MACRO sdffphc_2
  CLASS  CORE ;
  FOREIGN sdffphc_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 31.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 25.800 8.450 27.800 9.050 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 19.050 0.000 19.650 2.700 ;
        RECT 0.000 0.000 31.250 2.500 ;
        RECT 25.050 0.000 25.650 2.800 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.250 7.200 3.250 7.800 ;
    END
  END d
  PIN se
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.250 5.950 9.850 8.950 ;
        RECT 9.250 5.950 13.000 6.550 ;
        RECT 12.300 5.800 13.000 6.550 ;
    END
  END se
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 19.100 13.550 19.700 16.250 ;
        RECT 0.000 13.750 31.250 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 22.700 8.450 24.700 9.050 ;
    END
  END qb
  PIN g
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.750 7.200 6.400 7.800 ;
    END
  END g
  PIN sdi
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 11.250 9.700 13.250 10.300 ;
    END
  END sdi
  PIN clb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 9.700 2.250 10.300 ;
    END
  END clb
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 28.500 8.450 30.500 9.050 ;
    END
  END ck
  OBS 
      LAYER Metal1 ;
        RECT 1.450 8.450 8.350 9.050 ;
        RECT 10.550 7.550 13.750 8.150 ;
        RECT 10.550 7.550 11.150 9.050 ;
        RECT 15.950 5.800 16.550 6.550 ;
        RECT 14.250 5.950 16.550 6.550 ;
        RECT 14.250 5.950 14.850 9.200 ;
        RECT 14.250 8.600 17.050 9.200 ;
        RECT 17.250 5.950 21.350 6.550 ;
        RECT 17.250 5.950 17.850 7.650 ;
        RECT 15.350 7.050 17.850 7.650 ;
        RECT 15.350 7.050 15.950 8.100 ;
        RECT 7.000 4.700 22.700 5.300 ;
        RECT 22.100 4.700 22.700 6.700 ;
        RECT 22.100 6.100 25.250 6.700 ;
        RECT 19.450 7.200 30.850 7.800 ;
        RECT 19.450 7.200 20.050 8.750 ;
        RECT 17.550 8.150 20.050 8.750 ;
  END 
END sdffphc_2

MACRO sdffphc_1
  CLASS  CORE ;
  FOREIGN sdffphc_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 31.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 29.000 5.950 31.000 6.550 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 27.650 0.000 28.250 2.700 ;
        RECT 0.000 0.000 31.250 2.500 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.250 7.200 3.250 7.800 ;
    END
  END d
  PIN se
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.250 5.950 9.850 8.950 ;
        RECT 9.250 5.950 12.900 6.550 ;
        RECT 12.200 5.800 12.900 6.550 ;
    END
  END se
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 19.400 13.550 20.000 16.250 ;
        RECT 0.000 13.750 31.250 16.250 ;
        RECT 27.600 13.550 28.200 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 27.050 8.450 29.050 9.050 ;
    END
  END qb
  PIN g
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.750 7.200 6.400 7.800 ;
    END
  END g
  PIN sdi
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 12.000 9.700 14.000 10.300 ;
    END
  END sdi
  PIN clb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 9.700 2.250 10.300 ;
    END
  END clb
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 19.600 3.450 21.600 4.050 ;
    END
  END ck
  OBS 
      LAYER Metal1 ;
        RECT 1.450 8.450 8.350 9.050 ;
        RECT 10.550 7.550 13.750 8.150 ;
        RECT 10.550 7.550 11.150 9.050 ;
        RECT 15.850 5.800 16.450 7.000 ;
        RECT 14.250 6.400 16.450 7.000 ;
        RECT 14.250 6.400 14.850 9.200 ;
        RECT 14.250 8.600 17.050 9.200 ;
        RECT 17.000 5.950 23.150 6.550 ;
        RECT 17.000 5.950 17.600 8.100 ;
        RECT 15.350 7.500 17.600 8.100 ;
        RECT 22.550 8.450 25.750 9.050 ;
        RECT 18.100 7.200 26.450 7.800 ;
        RECT 18.100 7.200 18.700 7.950 ;
  END 
END sdffphc_1

MACRO sdffph_8
  CLASS  CORE ;
  FOREIGN sdffph_8 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 38.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 33.300 5.950 35.300 6.550 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 17.050 0.000 17.650 2.800 ;
        RECT 0.000 0.000 38.750 2.500 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.750 7.150 2.800 7.850 ;
    END
  END d
  PIN se
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.300 7.200 11.100 7.800 ;
    END
  END se
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 3.950 13.450 4.550 16.250 ;
        RECT 0.000 13.750 38.750 16.250 ;
        RECT 28.950 13.450 29.550 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 29.750 8.450 31.750 9.050 ;
    END
  END qb
  PIN g
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.400 7.200 5.400 7.800 ;
    END
  END g
  PIN sdi
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 10.850 4.700 12.850 5.300 ;
    END
  END sdi
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 36.150 4.700 38.200 5.300 ;
    END
  END ck
  OBS 
      LAYER Metal1 ;
        RECT 1.000 5.950 7.400 6.550 ;
        RECT 5.900 5.950 6.500 9.050 ;
        RECT 5.900 8.450 7.500 9.050 ;
        RECT 11.700 5.950 13.050 6.550 ;
        RECT 11.700 5.950 12.300 9.050 ;
        RECT 8.650 8.450 13.900 9.050 ;
        RECT 14.200 6.100 15.000 6.700 ;
        RECT 14.400 6.100 15.000 10.350 ;
        RECT 14.400 9.750 15.800 10.350 ;
        RECT 15.500 5.950 23.400 6.550 ;
        RECT 15.500 5.950 16.100 9.050 ;
        RECT 15.500 8.450 21.700 9.050 ;
        RECT 19.700 9.600 20.300 10.300 ;
        RECT 19.700 9.700 27.850 10.300 ;
        RECT 20.950 4.700 33.350 5.300 ;
        RECT 23.800 7.050 24.400 7.850 ;
        RECT 16.800 7.250 38.050 7.850 ;
  END 
END sdffph_8

MACRO sdffph_6
  CLASS  CORE ;
  FOREIGN sdffph_6 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 37.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 32.000 9.700 34.000 10.300 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 3.850 0.000 4.450 2.800 ;
        RECT 0.000 0.000 37.500 2.500 ;
        RECT 31.300 0.000 31.900 2.800 ;
        RECT 24.900 0.000 25.500 2.800 ;
        RECT 11.550 0.000 12.150 2.750 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.400 8.450 2.400 9.050 ;
    END
  END d
  PIN se
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.350 7.200 11.000 7.800 ;
    END
  END se
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 4.100 13.450 4.700 16.250 ;
        RECT 0.000 13.750 37.500 16.250 ;
        RECT 31.300 13.450 31.900 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 26.600 8.450 28.600 9.050 ;
    END
  END qb
  PIN g
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.900 7.200 5.600 7.800 ;
    END
  END g
  PIN sdi
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 10.900 4.700 12.900 5.300 ;
    END
  END sdi
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 35.000 5.950 37.000 6.550 ;
    END
  END ck
  OBS 
      LAYER Metal1 ;
        RECT 0.450 9.700 7.650 10.300 ;
        RECT 8.500 5.950 12.900 6.550 ;
        RECT 12.300 5.950 12.900 10.300 ;
        RECT 8.750 9.700 12.900 10.300 ;
        RECT 13.400 4.900 15.050 5.500 ;
        RECT 13.400 4.900 14.000 10.300 ;
        RECT 13.400 9.700 15.050 10.300 ;
        RECT 15.300 6.000 23.550 6.600 ;
        RECT 15.300 6.000 15.900 9.000 ;
        RECT 15.300 8.300 16.050 9.000 ;
        RECT 15.300 8.400 20.400 9.000 ;
        RECT 18.500 9.500 19.300 10.250 ;
        RECT 18.500 9.650 30.200 10.250 ;
        RECT 25.250 7.100 31.500 7.700 ;
        RECT 25.250 7.100 25.850 9.000 ;
        RECT 21.100 8.400 25.850 9.000 ;
        RECT 24.150 6.000 33.250 6.600 ;
        RECT 32.650 6.000 33.250 7.800 ;
        RECT 16.550 7.200 17.150 7.900 ;
        RECT 32.650 7.200 37.050 7.800 ;
        RECT 24.150 6.000 24.750 7.900 ;
        RECT 16.550 7.300 24.750 7.900 ;
  END 
END sdffph_6

MACRO sdffph_4
  CLASS  CORE ;
  FOREIGN sdffph_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 33.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 29.200 7.200 31.200 7.800 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 33.750 2.500 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.950 6.600 1.550 10.300 ;
        RECT 0.950 9.700 5.300 10.300 ;
        RECT 0.950 6.600 2.050 7.200 ;
    END
  END d
  PIN se
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.250 4.650 10.250 5.300 ;
    END
  END se
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 33.750 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 25.500 5.950 27.500 6.550 ;
    END
  END qb
  PIN g
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.350 4.700 0.950 5.900 ;
        RECT 0.350 4.700 1.950 5.300 ;
    END
  END g
  PIN sdi
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 10.900 4.700 11.500 7.800 ;
        RECT 10.900 4.700 11.550 5.300 ;
        RECT 9.900 7.200 11.500 7.800 ;
    END
  END sdi
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 16.700 5.950 18.700 6.550 ;
    END
  END ck
  OBS 
      LAYER Metal1 ;
        RECT 2.550 4.600 5.350 5.200 ;
        RECT 4.750 4.600 5.350 6.650 ;
        RECT 4.750 6.050 6.250 6.650 ;
        RECT 5.650 6.050 6.250 7.650 ;
        RECT 5.650 7.050 8.200 7.650 ;
        RECT 2.550 4.600 3.150 9.050 ;
        RECT 2.550 8.450 4.000 9.050 ;
        RECT 5.900 4.950 7.350 5.550 ;
        RECT 6.750 4.950 7.350 6.550 ;
        RECT 6.750 5.950 9.300 6.550 ;
        RECT 8.700 5.950 9.300 9.050 ;
        RECT 8.700 8.450 11.600 9.050 ;
        RECT 12.150 5.000 13.750 5.600 ;
        RECT 12.150 5.000 12.750 7.050 ;
        RECT 12.100 6.450 12.700 9.300 ;
        RECT 12.100 8.700 13.800 9.300 ;
        RECT 13.200 7.550 14.900 8.150 ;
        RECT 14.300 7.550 14.900 9.050 ;
        RECT 14.300 8.450 24.350 9.050 ;
        RECT 23.700 8.450 24.350 9.250 ;
        RECT 13.250 6.250 16.000 6.850 ;
        RECT 15.400 6.250 16.000 7.950 ;
        RECT 15.400 7.350 25.500 7.950 ;
        RECT 3.650 7.150 5.150 7.750 ;
        RECT 4.550 7.150 5.150 8.750 ;
        RECT 4.550 8.150 7.750 8.750 ;
        RECT 7.150 8.150 7.750 10.400 ;
        RECT 27.200 8.100 27.800 10.400 ;
        RECT 7.150 9.800 27.800 10.400 ;
  END 
END sdffph_4

MACRO sdffph_3
  CLASS  CORE ;
  FOREIGN sdffph_3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 31.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 27.500 5.950 29.500 6.550 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 31.250 2.500 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.650 6.600 1.250 10.300 ;
        RECT 0.650 9.700 5.350 10.300 ;
        RECT 0.650 6.600 2.050 7.200 ;
    END
  END d
  PIN se
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.600 4.700 10.600 5.300 ;
    END
  END se
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 16.600 13.550 17.200 16.250 ;
        RECT 0.000 13.750 31.250 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 24.300 5.950 26.300 6.550 ;
    END
  END qb
  PIN g
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.350 4.700 0.950 5.700 ;
        RECT 0.350 4.700 2.350 5.300 ;
    END
  END g
  PIN sdi
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 10.000 7.100 11.650 7.900 ;
    END
  END sdi
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 16.900 5.950 18.900 6.550 ;
    END
  END ck
  OBS 
      LAYER Metal1 ;
        RECT 3.100 5.950 6.150 6.550 ;
        RECT 5.550 5.950 6.150 7.900 ;
        RECT 5.550 7.300 8.400 7.900 ;
        RECT 3.100 5.950 3.700 9.050 ;
        RECT 6.100 4.850 7.650 5.450 ;
        RECT 7.050 4.850 7.650 6.550 ;
        RECT 7.050 5.950 9.500 6.550 ;
        RECT 8.900 5.950 9.500 9.050 ;
        RECT 8.900 8.450 11.800 9.050 ;
        RECT 12.250 4.900 13.950 5.500 ;
        RECT 12.250 4.900 12.850 7.950 ;
        RECT 12.300 7.350 12.900 9.300 ;
        RECT 12.300 8.700 14.000 9.300 ;
        RECT 13.400 7.550 15.100 8.150 ;
        RECT 14.500 7.550 15.100 9.050 ;
        RECT 14.500 8.450 24.400 9.050 ;
        RECT 13.350 6.200 16.200 6.800 ;
        RECT 15.600 6.200 16.200 7.950 ;
        RECT 15.600 7.350 24.400 7.950 ;
        RECT 4.200 7.300 4.800 9.000 ;
        RECT 4.200 8.400 6.500 9.000 ;
        RECT 5.900 8.400 6.500 10.400 ;
        RECT 15.850 9.550 27.000 10.150 ;
        RECT 26.400 7.350 27.000 10.150 ;
        RECT 5.900 9.800 16.450 10.400 ;
  END 
END sdffph_3

MACRO sdffph_2
  CLASS  CORE ;
  FOREIGN sdffph_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 28.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 23.400 8.400 25.300 9.100 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 3.350 0.000 3.950 2.650 ;
        RECT 0.000 0.000 28.750 2.500 ;
        RECT 22.550 0.000 23.150 2.800 ;
        RECT 16.550 0.000 17.150 2.700 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.500 8.400 2.300 9.100 ;
    END
  END d
  PIN se
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.050 7.500 6.650 9.050 ;
        RECT 6.050 7.500 7.900 8.100 ;
        RECT 5.950 8.350 6.650 9.050 ;
    END
  END se
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 3.450 13.550 4.050 16.250 ;
        RECT 0.000 13.750 28.750 16.250 ;
        RECT 16.600 13.550 17.200 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 20.700 8.450 22.700 9.050 ;
    END
  END qb
  PIN g
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.850 6.650 3.450 9.150 ;
        RECT 2.850 8.450 4.400 9.150 ;
    END
  END g
  PIN sdi
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.500 8.000 10.400 9.150 ;
        RECT 9.500 8.450 10.800 9.150 ;
    END
  END sdi
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 26.000 8.450 28.000 9.050 ;
    END
  END ck
  OBS 
      LAYER Metal1 ;
        RECT 6.050 5.800 8.650 6.400 ;
        RECT 9.750 5.650 10.350 7.500 ;
        RECT 8.400 6.900 11.500 7.500 ;
        RECT 10.900 6.900 11.500 7.950 ;
        RECT 8.400 6.900 9.000 9.200 ;
        RECT 7.900 8.600 9.000 9.200 ;
        RECT 13.450 5.800 14.050 6.550 ;
        RECT 12.000 5.950 14.050 6.550 ;
        RECT 12.000 5.950 12.600 9.200 ;
        RECT 12.000 8.600 14.500 9.200 ;
        RECT 14.850 6.250 18.850 6.850 ;
        RECT 14.850 6.250 15.450 7.650 ;
        RECT 13.150 7.050 15.450 7.650 ;
        RECT 13.150 7.050 13.750 8.100 ;
        RECT 8.650 4.550 11.450 5.150 ;
        RECT 4.900 4.700 9.250 5.300 ;
        RECT 10.850 4.700 20.200 5.300 ;
        RECT 19.600 4.700 20.200 6.750 ;
        RECT 19.600 6.150 22.750 6.750 ;
        RECT 4.900 4.700 5.500 7.800 ;
        RECT 19.550 7.250 28.350 7.850 ;
        RECT 16.950 7.350 20.150 7.950 ;
        RECT 16.950 7.350 17.550 8.750 ;
        RECT 15.000 8.150 17.550 8.750 ;
  END 
END sdffph_2

MACRO sdffph_1
  CLASS  CORE ;
  FOREIGN sdffph_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 28.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 26.500 5.950 28.500 6.550 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 3.350 0.000 3.950 2.700 ;
        RECT 0.000 0.000 28.750 2.500 ;
        RECT 25.150 0.000 25.750 2.700 ;
        RECT 6.200 0.000 6.800 2.700 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.800 8.450 2.800 9.050 ;
    END
  END d
  PIN se
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.850 7.200 7.900 7.850 ;
    END
  END se
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 3.450 13.550 4.050 16.250 ;
        RECT 0.000 13.750 28.750 16.250 ;
        RECT 25.100 13.550 25.700 16.250 ;
        RECT 16.900 13.550 17.500 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 25.000 8.450 27.000 9.050 ;
    END
  END qb
  PIN g
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.850 5.950 4.050 6.550 ;
        RECT 3.450 8.450 4.300 9.150 ;
        RECT 3.450 5.950 4.050 9.150 ;
    END
  END g
  PIN sdi
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.600 8.350 11.100 9.150 ;
    END
  END sdi
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 17.000 3.450 19.000 4.050 ;
    END
  END ck
  OBS 
      LAYER Metal1 ;
        RECT 0.350 3.450 6.650 4.050 ;
        RECT 6.050 5.950 8.750 6.550 ;
        RECT 10.600 5.300 12.150 5.900 ;
        RECT 10.600 5.300 11.200 6.600 ;
        RECT 9.850 6.000 11.200 6.600 ;
        RECT 9.850 6.000 10.450 7.800 ;
        RECT 8.450 7.200 10.450 7.800 ;
        RECT 8.450 7.200 9.050 9.200 ;
        RECT 7.900 8.600 9.050 9.200 ;
        RECT 13.350 5.800 13.950 7.000 ;
        RECT 11.750 6.400 13.950 7.000 ;
        RECT 11.750 6.400 12.350 9.200 ;
        RECT 11.750 8.600 14.550 9.200 ;
        RECT 14.500 6.250 20.650 6.850 ;
        RECT 14.500 6.250 15.100 8.100 ;
        RECT 12.850 7.500 15.100 8.100 ;
        RECT 20.050 8.450 23.250 9.050 ;
        RECT 15.600 7.350 23.950 7.950 ;
  END 
END sdffph_1

MACRO sdffpc_8
  CLASS  CORE ;
  FOREIGN sdffpc_8 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 35.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 29.350 8.450 31.350 9.050 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 35.000 2.500 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.450 4.700 3.350 5.800 ;
        RECT 2.450 4.700 4.450 5.300 ;
    END
  END d
  PIN se
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.500 8.450 5.750 9.100 ;
    END
  END se
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 7.100 13.450 7.700 16.250 ;
        RECT 0.000 13.750 35.000 16.250 ;
        RECT 25.100 13.450 25.700 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 25.900 8.450 27.900 9.050 ;
    END
  END qb
  PIN sdi
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.450 4.700 9.500 5.300 ;
    END
  END sdi
  PIN clb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.250 7.200 3.250 7.800 ;
    END
  END clb
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 32.300 4.700 34.350 5.300 ;
    END
  END ck
  OBS 
      LAYER Metal1 ;
        RECT 3.900 7.200 8.500 7.800 ;
        RECT 7.900 7.200 8.500 8.400 ;
        RECT 3.200 9.700 10.300 10.300 ;
        RECT 3.900 5.950 10.400 6.550 ;
        RECT 10.900 4.900 12.100 5.500 ;
        RECT 10.900 4.900 11.500 10.300 ;
        RECT 10.900 9.700 12.100 10.300 ;
        RECT 13.200 5.950 20.950 6.550 ;
        RECT 12.000 6.000 13.800 6.600 ;
        RECT 12.000 6.000 12.600 9.000 ;
        RECT 12.000 8.400 17.850 9.000 ;
        RECT 15.500 9.500 24.000 10.100 ;
        RECT 18.350 4.700 29.500 5.300 ;
        RECT 17.250 7.100 17.850 7.800 ;
        RECT 19.900 7.050 20.500 7.800 ;
        RECT 13.100 7.200 34.200 7.800 ;
        RECT 13.100 7.200 13.700 7.900 ;
  END 
END sdffpc_8

MACRO sdffpc_6
  CLASS  CORE ;
  FOREIGN sdffpc_6 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 33.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 28.250 9.700 30.350 10.300 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 27.550 0.000 28.150 2.650 ;
        RECT 0.000 0.000 33.750 2.500 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.200 4.700 2.800 5.900 ;
        RECT 2.200 4.700 4.050 5.300 ;
    END
  END d
  PIN se
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.500 8.450 2.850 9.050 ;
        RECT 2.250 8.700 5.300 9.300 ;
        RECT 4.700 8.450 5.300 9.300 ;
    END
  END se
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 6.400 13.450 7.000 16.250 ;
        RECT 0.000 13.750 33.750 16.250 ;
        RECT 27.550 13.450 28.150 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 22.850 8.450 24.850 9.050 ;
    END
  END qb
  PIN sdi
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.900 4.700 9.900 5.300 ;
    END
  END sdi
  PIN clb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.500 7.200 2.500 7.800 ;
    END
  END clb
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 31.250 5.950 33.250 6.550 ;
    END
  END ck
  OBS 
      LAYER Metal1 ;
        RECT 3.000 7.250 7.750 7.850 ;
        RECT 3.000 7.250 4.100 7.900 ;
        RECT 3.500 7.250 4.100 8.000 ;
        RECT 3.600 5.950 9.900 6.550 ;
        RECT 8.600 5.950 9.200 10.300 ;
        RECT 6.250 9.700 9.600 10.300 ;
        RECT 2.500 9.800 6.850 10.400 ;
        RECT 10.400 4.850 11.600 5.450 ;
        RECT 10.400 4.850 11.000 10.300 ;
        RECT 10.400 9.700 11.600 10.300 ;
        RECT 11.500 5.950 19.050 6.550 ;
        RECT 11.500 5.950 12.100 8.900 ;
        RECT 11.500 8.300 16.650 8.900 ;
        RECT 14.750 9.650 26.450 10.250 ;
        RECT 21.500 7.100 27.750 7.700 ;
        RECT 21.500 7.100 22.100 8.950 ;
        RECT 17.350 8.350 22.100 8.950 ;
        RECT 20.400 6.000 29.500 6.600 ;
        RECT 28.900 6.000 29.500 7.800 ;
        RECT 12.700 7.200 21.000 7.800 ;
        RECT 28.900 7.200 33.300 7.800 ;
        RECT 20.400 6.000 21.000 7.850 ;
        RECT 18.450 7.200 21.000 7.850 ;
  END 
END sdffpc_6

MACRO sdffpc_4
  CLASS  CORE ;
  FOREIGN sdffpc_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 30.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 25.550 7.200 27.550 7.800 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 30.000 2.500 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 8.350 2.200 9.050 ;
    END
  END d
  PIN se
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.750 3.450 5.750 4.050 ;
    END
  END se
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 30.000 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 21.750 5.950 23.850 6.550 ;
    END
  END qb
  PIN sdi
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.450 8.350 7.950 9.150 ;
    END
  END sdi
  PIN clb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.450 5.950 3.450 6.550 ;
    END
  END clb
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 13.450 5.950 14.750 6.550 ;
        RECT 14.150 5.950 14.750 8.200 ;
    END
  END ck
  OBS 
      LAYER Metal1 ;
        RECT 0.350 5.950 0.950 7.800 ;
        RECT 4.250 6.900 4.850 7.800 ;
        RECT 0.350 7.200 4.850 7.800 ;
        RECT 2.700 7.200 3.300 9.200 ;
        RECT 5.950 6.250 8.250 6.850 ;
        RECT 5.950 6.250 6.550 7.850 ;
        RECT 5.350 7.250 5.950 9.200 ;
        RECT 4.400 8.600 5.950 9.200 ;
        RECT 9.650 6.200 10.800 6.800 ;
        RECT 9.650 6.200 10.250 7.950 ;
        RECT 8.650 7.350 10.250 7.950 ;
        RECT 8.650 7.350 9.250 10.500 ;
        RECT 8.650 9.900 10.450 10.500 ;
        RECT 9.750 8.450 12.450 9.050 ;
        RECT 17.200 8.450 21.450 9.050 ;
        RECT 11.850 8.450 12.450 10.500 ;
        RECT 17.200 8.450 17.800 10.500 ;
        RECT 11.850 9.900 17.800 10.500 ;
        RECT 10.750 7.350 13.550 7.950 ;
        RECT 15.550 7.350 21.450 7.950 ;
        RECT 12.950 7.350 13.550 9.400 ;
        RECT 15.550 7.350 16.150 9.400 ;
        RECT 12.950 8.800 16.150 9.400 ;
  END 
END sdffpc_4

MACRO sdffpc_3
  CLASS  CORE ;
  FOREIGN sdffpc_3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 27.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 24.050 5.950 26.050 6.550 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 15.800 0.000 16.400 2.700 ;
        RECT 0.000 0.000 27.500 2.500 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 8.400 2.150 9.050 ;
    END
  END d
  PIN se
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.550 4.600 5.450 5.200 ;
        RECT 3.950 4.600 5.450 5.400 ;
    END
  END se
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 27.500 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 20.750 5.950 22.750 6.550 ;
    END
  END qb
  PIN sdi
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.450 8.450 8.450 9.050 ;
    END
  END sdi
  PIN clb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.950 4.650 2.850 5.350 ;
    END
  END clb
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 14.100 5.950 14.800 6.750 ;
        RECT 14.100 5.950 16.100 6.550 ;
    END
  END ck
  OBS 
      LAYER Metal1 ;
        RECT 0.350 5.950 1.000 7.800 ;
        RECT 3.950 6.900 4.550 7.800 ;
        RECT 0.350 7.200 4.550 7.800 ;
        RECT 2.700 7.200 3.300 9.200 ;
        RECT 5.650 6.900 6.250 7.850 ;
        RECT 5.050 7.250 8.450 7.850 ;
        RECT 5.050 7.250 5.650 9.200 ;
        RECT 4.400 8.600 5.650 9.200 ;
        RECT 8.950 5.950 10.650 6.550 ;
        RECT 8.950 5.950 9.550 10.200 ;
        RECT 8.950 9.600 10.900 10.200 ;
        RECT 10.050 8.450 20.650 9.050 ;
        RECT 10.500 7.150 11.100 7.950 ;
        RECT 10.500 7.350 20.650 7.950 ;
  END 
END sdffpc_3

MACRO sdffpc_2
  CLASS  CORE ;
  FOREIGN sdffpc_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 25.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 19.800 8.450 21.800 9.050 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 12.800 0.000 13.400 2.700 ;
        RECT 0.000 0.000 25.000 2.500 ;
        RECT 18.800 0.000 19.400 2.800 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 8.350 1.750 9.150 ;
    END
  END d
  PIN se
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.000 12.200 6.000 12.800 ;
    END
  END se
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 1.000 13.550 1.600 16.250 ;
        RECT 0.000 13.750 25.000 16.250 ;
        RECT 12.900 13.550 13.500 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 16.950 8.450 18.950 9.050 ;
    END
  END qb
  PIN sdi
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.650 8.350 7.150 9.150 ;
    END
  END sdi
  PIN clb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.450 5.850 2.950 6.650 ;
    END
  END clb
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 22.750 8.450 24.750 9.050 ;
    END
  END ck
  OBS 
      LAYER Metal1 ;
        RECT 3.450 6.150 4.650 6.750 ;
        RECT 0.350 5.950 0.950 7.800 ;
        RECT 3.450 6.150 4.050 7.800 ;
        RECT 0.350 7.200 4.050 7.800 ;
        RECT 2.700 7.200 3.300 9.200 ;
        RECT 6.550 5.300 8.350 5.900 ;
        RECT 6.550 5.300 7.150 6.750 ;
        RECT 5.750 6.150 7.150 6.750 ;
        RECT 5.750 6.150 6.350 7.850 ;
        RECT 4.550 7.250 6.350 7.850 ;
        RECT 4.550 7.250 5.150 9.200 ;
        RECT 4.400 8.600 5.150 9.200 ;
        RECT 9.050 5.800 10.300 6.400 ;
        RECT 7.950 6.400 9.650 7.000 ;
        RECT 7.950 6.400 8.550 9.200 ;
        RECT 7.950 8.600 10.750 9.200 ;
        RECT 11.000 6.250 15.100 6.850 ;
        RECT 10.150 7.050 11.600 7.650 ;
        RECT 11.000 6.250 11.600 7.650 ;
        RECT 9.050 7.500 10.750 8.100 ;
        RECT 15.800 7.250 24.600 7.850 ;
        RECT 13.200 7.350 16.400 7.950 ;
        RECT 13.200 7.350 13.800 8.750 ;
        RECT 11.250 8.150 13.800 8.750 ;
  END 
END sdffpc_2

MACRO sdffpc_1
  CLASS  CORE ;
  FOREIGN sdffpc_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 23.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 21.500 5.950 23.500 6.550 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 3.300 0.000 4.000 2.600 ;
        RECT 0.000 0.000 23.750 2.500 ;
        RECT 21.050 0.000 21.650 2.700 ;
        RECT 14.950 0.000 15.550 2.700 ;
        RECT 12.350 0.000 12.950 2.700 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 8.400 2.150 9.050 ;
    END
  END d
  PIN se
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.500 12.200 5.500 12.800 ;
    END
  END se
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 1.000 13.550 1.600 16.250 ;
        RECT 0.000 13.750 23.750 16.250 ;
        RECT 21.000 13.550 21.600 16.250 ;
        RECT 13.050 13.550 13.650 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 20.250 8.450 22.250 9.050 ;
    END
  END qb
  PIN sdi
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.650 8.350 7.150 9.150 ;
    END
  END sdi
  PIN clb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.450 5.850 2.950 6.650 ;
    END
  END clb
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 12.400 3.450 14.400 4.050 ;
    END
  END ck
  OBS 
      LAYER Metal1 ;
        RECT 3.450 6.150 4.650 6.750 ;
        RECT 0.350 5.950 0.950 7.800 ;
        RECT 3.450 6.150 4.050 7.800 ;
        RECT 0.350 7.200 4.050 7.800 ;
        RECT 2.700 7.200 3.300 9.200 ;
        RECT 6.550 5.300 8.150 5.900 ;
        RECT 6.550 5.300 7.150 6.750 ;
        RECT 5.750 6.150 7.150 6.750 ;
        RECT 5.750 6.150 6.350 7.850 ;
        RECT 4.550 7.250 6.350 7.850 ;
        RECT 4.550 7.250 5.150 9.200 ;
        RECT 4.400 8.600 5.150 9.200 ;
        RECT 9.250 5.800 9.850 7.000 ;
        RECT 7.650 6.400 9.850 7.000 ;
        RECT 7.650 6.400 8.250 9.200 ;
        RECT 7.650 8.600 10.450 9.200 ;
        RECT 10.500 5.950 16.550 6.550 ;
        RECT 10.500 5.950 11.100 8.100 ;
        RECT 8.750 7.500 11.100 8.100 ;
        RECT 15.950 8.450 19.050 9.050 ;
        RECT 11.600 7.200 19.850 7.800 ;
        RECT 11.600 7.200 12.200 8.000 ;
  END 
END sdffpc_1

MACRO sdffp_8
  CLASS  CORE ;
  FOREIGN sdffp_8 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 32.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 27.000 5.900 29.000 6.550 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 3.450 0.000 4.050 2.800 ;
        RECT 0.000 0.000 32.500 2.500 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.300 5.950 2.250 6.550 ;
        RECT 1.650 5.950 2.250 7.050 ;
    END
  END d
  PIN se
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.850 7.200 3.450 9.050 ;
        RECT 2.850 7.200 5.200 7.800 ;
        RECT 2.200 8.450 3.450 9.050 ;
    END
  END se
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 3.600 13.450 4.200 16.250 ;
        RECT 0.000 13.750 32.500 16.250 ;
        RECT 22.750 13.450 23.350 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 23.300 8.450 25.300 9.050 ;
    END
  END qb
  PIN sdi
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.050 8.450 6.050 9.050 ;
    END
  END sdi
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 29.950 4.700 32.000 5.300 ;
    END
  END ck
  OBS 
      LAYER Metal1 ;
        RECT 0.350 4.700 7.150 5.300 ;
        RECT 6.550 4.700 7.150 10.300 ;
        RECT 8.250 5.950 8.850 10.300 ;
        RECT 9.350 5.900 10.550 6.550 ;
        RECT 9.350 5.950 18.150 6.550 ;
        RECT 9.350 5.900 9.950 9.050 ;
        RECT 9.350 8.450 14.850 9.050 ;
        RECT 13.150 9.600 13.750 10.300 ;
        RECT 13.150 9.700 21.650 10.300 ;
        RECT 15.550 4.700 27.150 5.300 ;
        RECT 10.450 7.200 31.850 7.800 ;
        RECT 17.550 7.200 18.150 7.900 ;
  END 
END sdffp_8

MACRO sdffp_6
  CLASS  CORE ;
  FOREIGN sdffp_6 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 30.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 24.500 9.700 26.600 10.300 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 3.050 0.000 3.650 2.800 ;
        RECT 0.000 0.000 30.000 2.500 ;
        RECT 23.800 0.000 24.400 2.650 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.400 5.950 2.400 6.550 ;
    END
  END d
  PIN se
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.700 6.450 4.300 9.050 ;
        RECT 2.200 8.450 4.300 9.050 ;
    END
  END se
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 3.400 13.450 4.000 16.250 ;
        RECT 0.000 13.750 30.000 16.250 ;
        RECT 23.800 13.450 24.400 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 19.100 8.450 21.100 9.050 ;
    END
  END qb
  PIN sdi
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.350 4.700 6.350 5.300 ;
    END
  END sdi
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 27.500 5.950 29.500 6.550 ;
    END
  END ck
  OBS 
      LAYER Metal1 ;
        RECT 6.000 8.000 6.600 10.300 ;
        RECT 0.450 9.700 7.100 10.300 ;
        RECT 7.600 4.900 8.800 5.500 ;
        RECT 7.600 4.900 8.200 10.300 ;
        RECT 7.600 9.700 8.800 10.300 ;
        RECT 10.000 5.950 16.150 6.550 ;
        RECT 8.700 6.000 10.600 6.600 ;
        RECT 8.700 6.000 9.300 9.000 ;
        RECT 8.700 8.400 13.950 9.000 ;
        RECT 14.450 4.700 21.400 5.300 ;
        RECT 11.850 9.500 12.450 10.250 ;
        RECT 11.850 9.650 22.700 10.250 ;
        RECT 17.750 7.100 24.000 7.700 ;
        RECT 17.750 7.100 18.350 8.950 ;
        RECT 14.450 8.350 18.350 8.950 ;
        RECT 16.650 6.000 25.750 6.600 ;
        RECT 25.150 6.000 25.750 7.800 ;
        RECT 25.150 7.200 29.550 7.800 ;
        RECT 16.650 6.000 17.250 7.850 ;
        RECT 9.800 7.250 17.250 7.850 ;
        RECT 9.800 7.250 10.400 7.900 ;
  END 
END sdffp_6

MACRO sdffp_4
  CLASS  CORE ;
  FOREIGN sdffp_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 30.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 25.000 7.200 27.000 7.800 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 30.000 2.500 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.600 6.800 3.450 7.800 ;
        RECT 2.600 7.200 4.350 7.800 ;
    END
  END d
  PIN se
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.350 5.850 0.950 7.800 ;
        RECT 1.150 7.200 1.750 9.150 ;
        RECT 0.350 7.200 1.750 7.800 ;
    END
  END se
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 30.000 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 21.750 5.950 23.750 6.550 ;
    END
  END qb
  PIN sdi
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.950 7.100 6.550 9.150 ;
    END
  END sdi
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 12.500 5.950 14.500 6.550 ;
    END
  END ck
  OBS 
      LAYER Metal1 ;
        RECT 4.700 5.850 8.250 6.450 ;
        RECT 9.150 5.850 10.100 6.450 ;
        RECT 9.150 5.850 9.750 7.950 ;
        RECT 8.250 7.350 9.750 7.950 ;
        RECT 8.250 7.350 8.850 10.200 ;
        RECT 8.250 9.600 10.050 10.200 ;
        RECT 9.350 8.450 21.750 9.050 ;
        RECT 10.300 6.950 10.900 7.950 ;
        RECT 10.300 7.350 21.750 7.950 ;
  END 
END sdffp_4

MACRO sdffp_3
  CLASS  CORE ;
  FOREIGN sdffp_3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 27.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 23.550 5.950 25.550 6.550 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 27.500 2.500 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.450 6.600 4.050 7.800 ;
        RECT 3.050 7.200 4.550 7.800 ;
    END
  END d
  PIN se
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.350 5.800 1.550 6.450 ;
        RECT 0.950 6.000 2.800 6.600 ;
        RECT 0.950 5.800 1.550 7.800 ;
    END
  END se
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 27.500 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 20.750 5.950 22.750 6.550 ;
    END
  END qb
  PIN sdi
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.500 5.950 7.500 6.550 ;
    END
  END sdi
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 12.950 5.950 14.950 6.550 ;
    END
  END ck
  OBS 
      LAYER Metal1 ;
        RECT 4.100 8.550 7.900 9.150 ;
        RECT 8.400 6.050 10.100 6.650 ;
        RECT 8.400 6.050 9.000 10.150 ;
        RECT 8.400 9.550 10.050 10.150 ;
        RECT 10.150 7.150 10.800 7.950 ;
        RECT 10.150 7.350 20.000 7.950 ;
        RECT 9.500 8.450 20.150 9.050 ;
        RECT 19.550 8.450 20.150 9.450 ;
  END 
END sdffp_3

MACRO sdffnr_8
  CLASS  CORE ;
  FOREIGN sdffnr_8 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 35.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 23.600 9.700 27.600 10.300 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 22.300 0.000 22.900 2.800 ;
        RECT 0.000 0.000 35.000 2.500 ;
        RECT 25.300 0.000 25.900 2.800 ;
    END
  END vss!
  PIN ckb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 32.500 4.700 34.500 5.300 ;
    END
  END ckb
  PIN se
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.150 7.250 4.750 9.050 ;
        RECT 4.150 7.250 7.300 7.850 ;
        RECT 1.600 8.350 4.750 9.050 ;
    END
  END se
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.800 4.700 7.400 6.650 ;
        RECT 6.800 4.700 7.800 5.300 ;
        RECT 4.850 5.850 7.400 6.650 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 1.700 13.500 2.300 16.250 ;
        RECT 0.000 13.750 35.000 16.250 ;
        RECT 32.100 13.450 32.700 16.250 ;
        RECT 25.300 13.450 25.900 16.250 ;
        RECT 20.550 13.450 21.150 16.250 ;
        RECT 4.800 13.450 5.400 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 29.550 8.450 31.550 9.050 ;
    END
  END qb
  PIN sdi
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.400 8.450 7.400 9.050 ;
        RECT 6.550 8.450 7.400 9.250 ;
    END
  END sdi
  PIN rb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.350 4.550 1.950 5.400 ;
    END
  END rb
  OBS 
      LAYER Metal1 ;
        RECT 2.450 4.650 6.300 5.250 ;
        RECT 2.450 4.650 3.050 7.650 ;
        RECT 1.600 7.050 3.050 7.650 ;
        RECT 0.400 5.900 1.650 6.500 ;
        RECT 7.900 6.200 9.500 6.800 ;
        RECT 0.400 9.700 1.600 10.300 ;
        RECT 0.400 5.900 1.000 10.300 ;
        RECT 7.900 6.200 8.500 10.400 ;
        RECT 1.000 9.800 8.500 10.400 ;
        RECT 10.100 5.150 11.200 5.750 ;
        RECT 10.100 5.150 10.700 7.950 ;
        RECT 9.000 7.350 10.700 7.950 ;
        RECT 9.000 7.350 9.600 10.300 ;
        RECT 9.000 9.700 10.700 10.300 ;
        RECT 16.250 7.150 16.900 7.950 ;
        RECT 12.400 7.350 16.900 7.950 ;
        RECT 13.650 4.600 21.650 5.200 ;
        RECT 13.650 4.600 14.250 5.750 ;
        RECT 21.050 4.600 21.650 6.800 ;
        RECT 14.400 9.650 22.850 10.250 ;
        RECT 17.550 6.800 18.150 9.150 ;
        RECT 22.250 8.450 26.250 9.050 ;
        RECT 17.550 8.550 22.850 9.150 ;
        RECT 24.000 5.300 29.700 5.900 ;
        RECT 15.150 5.700 19.350 6.300 ;
        RECT 18.750 5.700 19.350 6.950 ;
        RECT 11.300 6.250 15.750 6.850 ;
        RECT 18.750 6.350 20.550 6.950 ;
        RECT 19.950 6.350 20.550 7.950 ;
        RECT 28.050 7.200 34.400 7.800 ;
        RECT 19.950 7.350 28.650 7.950 ;
        RECT 11.300 6.250 11.900 9.050 ;
        RECT 10.100 8.450 15.950 9.050 ;
        RECT 15.350 8.450 15.950 9.100 ;
  END 
END sdffnr_8

MACRO sdffnr_6
  CLASS  CORE ;
  FOREIGN sdffnr_6 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 33.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 25.150 9.700 29.150 10.300 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 23.950 0.000 24.550 2.650 ;
        RECT 0.000 0.000 33.750 2.500 ;
        RECT 26.850 0.000 27.450 2.650 ;
        RECT 25.400 0.000 26.000 2.650 ;
    END
  END vss!
  PIN ckb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 32.900 6.050 33.500 10.300 ;
        RECT 32.200 9.700 33.500 10.300 ;
    END
  END ckb
  PIN se
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.650 4.650 5.650 5.300 ;
    END
  END se
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.650 4.700 2.250 5.500 ;
        RECT 0.850 4.700 2.850 5.400 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 33.750 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 20.450 9.700 24.450 10.300 ;
    END
  END qb
  PIN sdi
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.650 8.400 7.300 10.300 ;
        RECT 5.950 9.700 7.300 10.300 ;
    END
  END sdi
  PIN rb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.950 7.300 1.650 9.050 ;
        RECT 0.950 7.300 2.900 7.900 ;
        RECT 0.250 8.450 1.650 9.050 ;
    END
  END rb
  OBS 
      LAYER Metal1 ;
        RECT 0.350 6.000 4.050 6.600 ;
        RECT 3.450 7.300 5.000 7.900 ;
        RECT 3.450 6.000 4.050 9.250 ;
        RECT 2.700 8.650 4.050 9.250 ;
        RECT 5.550 7.300 9.150 7.900 ;
        RECT 5.550 7.300 6.150 9.000 ;
        RECT 4.600 8.400 6.150 9.000 ;
        RECT 4.600 8.400 5.200 9.600 ;
        RECT 10.600 5.700 11.200 6.500 ;
        RECT 16.300 5.850 17.250 6.500 ;
        RECT 9.650 5.900 17.250 6.500 ;
        RECT 9.650 5.900 10.250 10.300 ;
        RECT 9.650 9.700 11.850 10.300 ;
        RECT 26.850 7.900 30.850 8.700 ;
        RECT 30.250 7.900 30.850 9.800 ;
        RECT 20.350 6.450 31.000 7.050 ;
        RECT 10.750 8.100 14.750 8.700 ;
        RECT 20.350 6.450 20.950 9.050 ;
        RECT 18.450 8.450 20.950 9.050 ;
        RECT 14.150 8.100 14.750 10.300 ;
        RECT 18.450 8.450 19.050 10.300 ;
        RECT 14.150 9.650 19.050 10.300 ;
        RECT 19.050 4.750 32.600 5.350 ;
        RECT 11.650 7.000 16.700 7.600 ;
        RECT 19.050 4.750 19.650 7.950 ;
        RECT 15.950 7.350 19.650 7.950 ;
        RECT 31.800 4.750 32.400 8.000 ;
        RECT 15.950 7.000 16.550 9.150 ;
  END 
END sdffnr_6

MACRO sdffnr_4
  CLASS  CORE ;
  FOREIGN sdffnr_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 28.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 22.300 9.700 24.300 10.300 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 28.750 2.500 ;
    END
  END vss!
  PIN ckb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 27.900 5.900 28.500 10.300 ;
        RECT 27.200 9.700 28.500 10.300 ;
    END
  END ckb
  PIN se
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.650 4.600 5.750 5.300 ;
    END
  END se
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.650 4.700 2.250 5.450 ;
        RECT 1.000 4.700 2.850 5.400 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 28.750 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 19.300 9.700 21.300 10.300 ;
    END
  END qb
  PIN sdi
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.650 8.400 7.300 10.300 ;
        RECT 5.850 9.700 7.300 10.300 ;
    END
  END sdi
  PIN rb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.950 7.300 1.650 9.150 ;
        RECT 0.950 7.300 2.900 7.900 ;
        RECT 0.250 8.450 1.650 9.150 ;
    END
  END rb
  OBS 
      LAYER Metal1 ;
        RECT 0.350 6.000 4.050 6.600 ;
        RECT 3.450 7.300 5.000 7.900 ;
        RECT 3.450 6.000 4.050 9.250 ;
        RECT 2.700 8.650 4.050 9.250 ;
        RECT 5.550 7.300 9.150 7.900 ;
        RECT 5.550 7.300 6.150 9.000 ;
        RECT 4.600 8.400 6.150 9.000 ;
        RECT 4.600 8.400 5.200 9.600 ;
        RECT 16.350 5.850 16.950 6.500 ;
        RECT 9.650 5.900 16.950 6.500 ;
        RECT 9.650 5.900 10.250 10.300 ;
        RECT 9.650 9.700 11.350 10.300 ;
        RECT 20.050 6.450 26.000 7.050 ;
        RECT 20.050 6.450 20.650 9.050 ;
        RECT 18.150 8.450 20.650 9.050 ;
        RECT 10.750 8.600 14.300 9.200 ;
        RECT 13.700 8.450 14.300 10.200 ;
        RECT 18.150 8.450 18.750 10.200 ;
        RECT 13.700 9.550 18.750 10.200 ;
        RECT 18.550 4.700 27.550 5.300 ;
        RECT 10.800 7.200 11.400 7.950 ;
        RECT 26.800 4.700 27.400 7.800 ;
        RECT 18.550 4.700 19.150 7.950 ;
        RECT 10.800 7.350 19.150 7.950 ;
        RECT 15.600 7.350 16.200 9.050 ;
  END 
END sdffnr_4

MACRO sdffnr_3
  CLASS  CORE ;
  FOREIGN sdffnr_3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 27.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 21.550 9.700 23.550 10.300 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 27.500 2.500 ;
    END
  END vss!
  PIN ckb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 25.950 4.700 27.250 5.300 ;
        RECT 26.650 4.700 27.250 8.350 ;
    END
  END ckb
  PIN se
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.350 8.100 3.950 8.750 ;
        RECT 4.000 9.700 5.300 10.300 ;
        RECT 4.000 8.150 4.600 10.300 ;
        RECT 3.350 8.150 4.600 8.750 ;
    END
  END se
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.150 4.700 1.750 6.000 ;
        RECT 1.150 4.700 2.800 5.400 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 27.500 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 18.900 9.700 20.900 10.300 ;
    END
  END qb
  PIN sdi
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.700 8.400 7.350 10.300 ;
        RECT 6.700 9.700 7.950 10.300 ;
    END
  END sdi
  PIN rb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.450 7.650 1.050 9.050 ;
        RECT 0.450 8.450 1.700 9.050 ;
    END
  END rb
  OBS 
      LAYER Metal1 ;
        RECT 2.450 5.900 6.850 6.550 ;
        RECT 2.450 5.900 3.050 7.400 ;
        RECT 2.200 6.800 2.800 10.400 ;
        RECT 2.200 9.800 3.300 10.400 ;
        RECT 4.550 7.050 8.550 7.650 ;
        RECT 9.050 4.900 16.350 5.500 ;
        RECT 15.750 4.900 16.350 5.600 ;
        RECT 9.050 4.900 9.650 10.350 ;
        RECT 9.050 9.750 10.950 10.350 ;
        RECT 10.150 8.450 10.750 9.200 ;
        RECT 17.600 8.150 24.750 8.800 ;
        RECT 13.400 7.500 14.050 9.200 ;
        RECT 10.150 8.600 14.050 9.200 ;
        RECT 13.400 7.500 14.000 10.350 ;
        RECT 17.600 8.150 18.200 10.350 ;
        RECT 13.400 9.750 18.200 10.350 ;
        RECT 10.700 6.350 15.950 6.950 ;
        RECT 15.350 6.450 26.150 7.050 ;
        RECT 10.700 6.350 11.300 7.900 ;
        RECT 15.350 6.350 15.950 9.200 ;
        RECT 25.550 6.450 26.150 9.900 ;
        RECT 25.550 9.300 26.300 9.900 ;
  END 
END sdffnr_3

MACRO sdffp_2
  CLASS  CORE ;
  FOREIGN sdffp_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 23.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 18.550 8.450 20.550 9.050 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 3.350 0.000 3.950 2.650 ;
        RECT 0.000 0.000 23.750 2.500 ;
        RECT 17.550 0.000 18.150 2.800 ;
        RECT 11.550 0.000 12.150 2.700 ;
        RECT 4.450 0.000 5.050 2.650 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.900 5.950 5.500 6.950 ;
        RECT 4.300 5.950 5.800 6.650 ;
    END
  END d
  PIN se
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.950 6.500 3.550 9.100 ;
        RECT 2.950 8.400 4.250 9.100 ;
    END
  END se
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 3.450 13.550 4.050 16.250 ;
        RECT 0.000 13.750 23.750 16.250 ;
        RECT 11.600 13.550 12.200 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 15.200 8.450 17.200 9.050 ;
    END
  END qb
  PIN sdi
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.300 8.450 2.300 9.050 ;
    END
  END sdi
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 21.300 8.450 23.300 9.050 ;
    END
  END ck
  OBS 
      LAYER Metal1 ;
        RECT 8.450 5.800 9.050 6.550 ;
        RECT 6.400 5.950 9.050 6.550 ;
        RECT 6.400 5.950 7.000 9.200 ;
        RECT 6.400 8.600 9.200 9.200 ;
        RECT 9.750 5.950 13.850 6.550 ;
        RECT 9.750 5.950 10.350 7.650 ;
        RECT 7.500 7.050 10.350 7.650 ;
        RECT 7.500 7.050 8.100 8.100 ;
        RECT 11.950 7.200 23.350 7.800 ;
        RECT 11.950 7.200 12.550 8.750 ;
        RECT 10.000 8.150 12.550 8.750 ;
  END 
END sdffp_2

MACRO sdffp_1
  CLASS  CORE ;
  FOREIGN sdffp_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 22.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 20.250 5.950 22.250 6.550 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 3.350 0.000 3.950 2.650 ;
        RECT 0.000 0.000 22.500 2.500 ;
        RECT 19.800 0.000 20.400 2.700 ;
        RECT 13.700 0.000 14.300 2.700 ;
        RECT 11.100 0.000 11.700 2.700 ;
        RECT 4.450 0.000 5.050 2.650 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.900 5.950 5.500 7.150 ;
        RECT 4.050 5.950 5.900 6.550 ;
    END
  END d
  PIN se
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.950 6.700 3.550 9.200 ;
        RECT 2.950 8.450 4.250 9.200 ;
    END
  END se
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 3.450 13.550 4.050 16.250 ;
        RECT 0.000 13.750 22.500 16.250 ;
        RECT 19.750 13.550 20.350 16.250 ;
        RECT 11.550 13.550 12.150 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 19.000 8.450 21.000 9.050 ;
    END
  END qb
  PIN sdi
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.300 8.450 2.300 9.050 ;
    END
  END sdi
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 11.550 3.450 13.550 4.050 ;
    END
  END ck
  OBS 
      LAYER Metal1 ;
        RECT 8.000 5.800 8.600 6.550 ;
        RECT 6.400 5.950 8.600 6.550 ;
        RECT 6.400 5.950 7.000 9.200 ;
        RECT 6.400 8.600 9.200 9.200 ;
        RECT 9.250 5.950 15.300 6.550 ;
        RECT 9.250 5.950 9.850 8.100 ;
        RECT 7.500 7.500 9.850 8.100 ;
        RECT 14.700 8.450 17.900 9.050 ;
        RECT 10.350 7.200 18.600 7.800 ;
        RECT 10.350 7.200 10.950 7.950 ;
  END 
END sdffp_1

MACRO sdffnr_2
  CLASS  CORE ;
  FOREIGN sdffnr_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 26.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 20.750 9.700 22.750 10.300 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 11.050 0.000 11.650 2.700 ;
        RECT 0.000 0.000 26.250 2.500 ;
    END
  END vss!
  PIN ckb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 24.700 5.950 26.000 6.550 ;
        RECT 25.400 5.950 26.000 8.950 ;
    END
  END ckb
  PIN se
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.050 4.650 5.300 5.250 ;
        RECT 4.700 4.650 5.300 5.300 ;
    END
  END se
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.100 5.850 3.450 6.750 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 1.000 13.400 1.600 16.250 ;
        RECT 0.000 13.750 26.250 16.250 ;
        RECT 19.750 13.450 20.350 16.250 ;
        RECT 10.150 13.400 10.750 16.250 ;
        RECT 7.000 13.550 7.600 16.250 ;
        RECT 2.700 13.450 3.300 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 18.050 9.700 20.100 10.300 ;
    END
  END qb
  PIN sdi
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.200 8.350 7.900 9.150 ;
    END
  END sdi
  PIN rb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 8.350 1.750 9.150 ;
    END
  END rb
  OBS 
      LAYER Metal1 ;
        RECT 1.000 5.850 1.600 7.850 ;
        RECT 3.950 6.900 4.550 7.850 ;
        RECT 1.000 7.250 4.550 7.850 ;
        RECT 2.400 7.250 3.000 9.200 ;
        RECT 5.650 6.900 6.250 7.850 ;
        RECT 5.050 7.250 7.950 7.850 ;
        RECT 5.050 7.250 5.650 9.200 ;
        RECT 4.100 8.600 5.650 9.200 ;
        RECT 9.550 7.150 10.150 7.950 ;
        RECT 14.700 6.050 15.300 7.950 ;
        RECT 9.550 7.350 15.300 7.950 ;
        RECT 9.450 4.750 15.350 5.350 ;
        RECT 9.450 4.750 10.050 6.550 ;
        RECT 8.450 5.950 10.050 6.550 ;
        RECT 8.450 5.950 9.050 10.300 ;
        RECT 8.450 9.700 11.150 10.300 ;
        RECT 15.850 4.700 16.500 5.300 ;
        RECT 15.850 4.700 16.450 9.200 ;
        RECT 10.300 8.450 14.450 9.050 ;
        RECT 16.950 8.450 23.800 9.050 ;
        RECT 10.300 8.450 11.050 9.100 ;
        RECT 13.850 8.450 14.450 10.300 ;
        RECT 16.950 7.450 17.550 10.300 ;
        RECT 13.850 9.700 17.550 10.300 ;
        RECT 16.950 6.050 18.700 6.650 ;
        RECT 18.100 6.050 18.700 7.850 ;
        RECT 18.100 7.250 24.900 7.850 ;
        RECT 24.300 7.250 24.900 10.150 ;
  END 
END sdffnr_2

MACRO sdffnr_1
  CLASS  CORE ;
  FOREIGN sdffnr_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 26.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 20.750 5.950 22.750 6.550 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 11.100 0.000 11.700 2.700 ;
        RECT 0.000 0.000 26.250 2.500 ;
    END
  END vss!
  PIN ckb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 23.400 5.950 26.000 6.550 ;
        RECT 25.400 5.950 26.000 9.100 ;
    END
  END ckb
  PIN se
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.450 3.400 4.500 4.050 ;
    END
  END se
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.100 5.850 3.450 6.750 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 1.000 13.400 1.600 16.250 ;
        RECT 0.000 13.750 26.250 16.250 ;
        RECT 10.150 13.400 10.750 16.250 ;
        RECT 7.000 13.550 7.600 16.250 ;
        RECT 2.700 13.450 3.300 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 17.450 5.950 19.450 6.550 ;
    END
  END qb
  PIN sdi
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.150 8.350 7.950 9.100 ;
    END
  END sdi
  PIN rb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 8.350 1.900 9.100 ;
    END
  END rb
  OBS 
      LAYER Metal1 ;
        RECT 1.000 5.850 1.600 7.850 ;
        RECT 3.950 6.800 4.550 7.850 ;
        RECT 1.000 7.250 4.550 7.850 ;
        RECT 2.400 7.250 3.000 9.100 ;
        RECT 5.650 6.800 6.250 7.850 ;
        RECT 5.050 7.250 7.950 7.850 ;
        RECT 5.050 7.250 5.650 9.100 ;
        RECT 4.100 8.500 5.650 9.100 ;
        RECT 9.650 7.300 15.200 7.900 ;
        RECT 8.450 6.100 15.300 6.700 ;
        RECT 8.450 6.100 9.050 10.300 ;
        RECT 8.450 9.700 11.150 10.300 ;
        RECT 15.850 5.900 16.450 9.200 ;
        RECT 10.650 8.400 11.250 9.050 ;
        RECT 16.950 8.300 17.600 9.050 ;
        RECT 10.650 8.450 13.950 9.050 ;
        RECT 16.950 8.450 23.800 9.050 ;
        RECT 13.350 8.450 13.950 10.300 ;
        RECT 16.950 8.300 17.550 10.300 ;
        RECT 13.350 9.700 17.550 10.300 ;
        RECT 16.950 7.200 24.900 7.800 ;
        RECT 24.300 7.200 24.900 10.300 ;
  END 
END sdffnr_1

MACRO sdffnh_8
  CLASS  CORE ;
  FOREIGN sdffnh_8 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 37.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 32.000 8.450 34.000 9.050 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 16.850 0.000 17.450 2.800 ;
        RECT 0.000 0.000 37.500 2.500 ;
    END
  END vss!
  PIN ckb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 34.950 4.700 37.100 5.300 ;
    END
  END ckb
  PIN se
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.650 7.100 9.050 7.700 ;
        RECT 8.500 7.200 11.300 7.800 ;
    END
  END se
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.750 7.200 2.900 7.800 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 3.950 13.450 4.550 16.250 ;
        RECT 0.000 13.750 37.500 16.250 ;
        RECT 27.750 13.450 28.350 16.250 ;
        RECT 14.400 13.450 15.000 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 28.300 8.450 30.300 9.050 ;
    END
  END qb
  PIN g
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.400 7.200 5.400 7.800 ;
    END
  END g
  PIN sdi
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 10.700 4.700 12.700 5.300 ;
    END
  END sdi
  OBS 
      LAYER Metal1 ;
        RECT 5.900 5.800 7.150 6.400 ;
        RECT 1.000 5.950 6.500 6.550 ;
        RECT 5.900 5.800 6.500 8.800 ;
        RECT 5.900 8.200 7.650 8.800 ;
        RECT 8.750 8.600 13.250 9.200 ;
        RECT 14.300 5.800 14.900 7.950 ;
        RECT 14.750 7.350 15.350 9.200 ;
        RECT 22.650 7.050 23.250 7.800 ;
        RECT 16.950 7.200 23.250 7.800 ;
        RECT 16.950 7.200 17.550 7.950 ;
        RECT 24.750 7.050 25.350 9.050 ;
        RECT 21.750 8.450 25.350 9.050 ;
        RECT 5.750 9.300 6.350 10.300 ;
        RECT 19.650 9.600 20.250 10.300 ;
        RECT 5.750 9.700 26.650 10.300 ;
        RECT 20.850 4.700 32.150 5.300 ;
        RECT 15.400 5.950 36.850 6.550 ;
        RECT 15.850 5.950 16.450 9.050 ;
        RECT 15.850 8.450 21.150 9.050 ;
  END 
END sdffnh_8

MACRO sdffnh_6
  CLASS  CORE ;
  FOREIGN sdffnh_6 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 36.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 30.750 9.700 32.850 10.300 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 3.850 0.000 4.450 2.800 ;
        RECT 0.000 0.000 36.250 2.500 ;
        RECT 30.050 0.000 30.650 2.800 ;
        RECT 23.650 0.000 24.250 2.800 ;
        RECT 11.550 0.000 12.150 2.800 ;
    END
  END vss!
  PIN ckb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 33.750 7.200 35.750 7.800 ;
    END
  END ckb
  PIN se
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.400 7.200 11.000 7.800 ;
    END
  END se
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.950 8.450 2.950 9.050 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 4.100 13.450 4.700 16.250 ;
        RECT 0.000 13.750 36.250 16.250 ;
        RECT 30.050 13.450 30.650 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 25.350 8.450 27.350 9.050 ;
    END
  END qb
  PIN g
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.100 7.200 5.600 7.800 ;
    END
  END g
  PIN sdi
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 10.500 4.700 12.500 5.300 ;
    END
  END sdi
  OBS 
      LAYER Metal1 ;
        RECT 0.700 9.700 7.650 10.300 ;
        RECT 8.500 5.950 13.000 6.550 ;
        RECT 12.400 5.950 13.000 10.300 ;
        RECT 8.750 9.700 13.000 10.300 ;
        RECT 14.000 5.200 14.700 5.800 ;
        RECT 14.000 5.200 14.600 10.300 ;
        RECT 14.000 9.650 15.050 10.300 ;
        RECT 16.300 7.200 19.900 7.800 ;
        RECT 18.100 9.500 18.700 10.250 ;
        RECT 18.100 9.650 28.950 10.250 ;
        RECT 24.000 7.100 30.250 7.700 ;
        RECT 24.000 7.100 24.600 9.150 ;
        RECT 20.700 8.550 24.600 9.150 ;
        RECT 20.700 4.850 33.650 5.450 ;
        RECT 15.200 5.950 22.450 6.550 ;
        RECT 21.850 6.000 35.800 6.600 ;
        RECT 15.200 8.300 20.000 8.900 ;
        RECT 15.200 5.950 15.800 9.000 ;
        RECT 15.100 8.400 15.800 9.000 ;
  END 
END sdffnh_6

MACRO sdffnh_4
  CLASS  CORE ;
  FOREIGN sdffnh_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 33.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 29.200 7.200 31.200 7.800 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 33.750 2.500 ;
    END
  END vss!
  PIN ckb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 16.900 5.950 18.900 6.550 ;
    END
  END ckb
  PIN se
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.450 4.700 10.500 5.300 ;
    END
  END se
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.950 6.350 1.550 10.300 ;
        RECT 0.950 9.700 5.100 10.300 ;
        RECT 4.150 9.450 5.100 10.300 ;
        RECT 0.950 6.350 2.100 7.100 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 20.350 13.450 21.050 16.250 ;
        RECT 0.000 13.750 33.750 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 25.500 5.950 27.500 6.550 ;
    END
  END qb
  PIN g
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.300 4.700 2.300 5.300 ;
    END
  END g
  PIN sdi
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 10.950 5.950 11.550 7.800 ;
        RECT 9.900 7.200 11.550 7.800 ;
    END
  END sdi
  OBS 
      LAYER Metal1 ;
        RECT 2.600 6.200 6.650 6.800 ;
        RECT 6.050 6.200 6.650 7.650 ;
        RECT 6.050 7.050 7.450 7.650 ;
        RECT 2.600 6.200 3.200 9.050 ;
        RECT 6.850 7.050 7.450 9.050 ;
        RECT 2.600 8.450 3.800 9.050 ;
        RECT 6.850 8.450 8.200 9.050 ;
        RECT 5.900 5.100 7.750 5.700 ;
        RECT 7.150 5.100 7.750 6.550 ;
        RECT 7.150 5.950 9.300 6.550 ;
        RECT 8.700 5.950 9.300 9.050 ;
        RECT 8.700 8.450 11.600 9.050 ;
        RECT 12.200 5.150 13.800 5.750 ;
        RECT 12.200 5.150 12.800 7.950 ;
        RECT 12.100 7.350 12.700 9.300 ;
        RECT 12.100 8.700 13.800 9.300 ;
        RECT 13.300 7.550 15.200 8.150 ;
        RECT 14.600 7.550 15.200 9.050 ;
        RECT 14.600 8.450 21.450 9.050 ;
        RECT 13.300 6.250 16.300 6.850 ;
        RECT 20.300 6.700 23.700 7.300 ;
        RECT 15.700 6.250 16.300 7.950 ;
        RECT 20.300 6.700 20.900 7.950 ;
        RECT 15.700 7.350 20.900 7.950 ;
        RECT 24.100 5.400 24.850 6.000 ;
        RECT 24.250 5.400 24.850 9.300 ;
        RECT 23.700 8.700 24.850 9.300 ;
        RECT 4.050 7.350 5.550 7.950 ;
        RECT 4.950 7.350 5.550 8.750 ;
        RECT 4.950 8.150 6.300 8.750 ;
        RECT 5.700 8.150 6.300 10.400 ;
        RECT 27.250 8.050 27.850 10.400 ;
        RECT 5.700 9.800 27.850 10.400 ;
  END 
END sdffnh_4

MACRO sdffnh_3
  CLASS  CORE ;
  FOREIGN sdffnh_3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 31.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 27.500 5.950 29.500 6.550 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 31.250 2.500 ;
    END
  END vss!
  PIN ckb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 16.900 5.950 18.900 6.550 ;
    END
  END ckb
  PIN se
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.100 4.700 11.100 5.300 ;
    END
  END se
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.950 6.400 1.550 10.300 ;
        RECT 0.950 9.700 5.150 10.300 ;
        RECT 4.150 9.250 5.150 10.300 ;
        RECT 0.950 6.400 2.050 7.100 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 31.250 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 24.600 5.950 26.600 6.550 ;
    END
  END qb
  PIN g
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.350 4.700 2.350 5.300 ;
    END
  END g
  PIN sdi
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 10.000 7.100 11.800 7.900 ;
    END
  END sdi
  OBS 
      LAYER Metal1 ;
        RECT 3.450 5.700 4.050 6.550 ;
        RECT 3.450 5.850 7.300 6.550 ;
        RECT 6.700 5.850 7.300 7.650 ;
        RECT 7.050 7.050 7.650 9.050 ;
        RECT 3.100 5.950 3.700 8.950 ;
        RECT 7.050 8.450 8.400 9.050 ;
        RECT 6.100 4.750 8.600 5.350 ;
        RECT 8.000 4.750 8.600 6.550 ;
        RECT 8.000 5.950 9.500 6.550 ;
        RECT 8.900 5.950 9.500 9.050 ;
        RECT 8.900 8.450 11.800 9.050 ;
        RECT 12.300 5.200 14.000 5.800 ;
        RECT 12.300 5.200 12.900 9.300 ;
        RECT 12.300 8.700 14.000 9.300 ;
        RECT 13.400 7.600 15.100 8.200 ;
        RECT 14.500 7.600 15.100 9.050 ;
        RECT 14.500 8.450 21.400 9.050 ;
        RECT 20.250 6.200 22.850 6.800 ;
        RECT 13.400 6.300 16.200 6.900 ;
        RECT 15.600 6.300 16.200 7.950 ;
        RECT 20.250 6.200 20.850 7.950 ;
        RECT 15.600 7.350 20.850 7.950 ;
        RECT 23.250 4.850 24.050 5.450 ;
        RECT 23.450 4.850 24.050 9.050 ;
        RECT 22.900 8.450 24.050 9.050 ;
        RECT 4.200 7.100 6.200 7.700 ;
        RECT 5.600 7.100 6.200 8.750 ;
        RECT 5.900 8.150 6.500 10.400 ;
        RECT 26.400 7.350 27.000 10.400 ;
        RECT 5.900 9.800 27.000 10.400 ;
  END 
END sdffnh_3

MACRO sdffnh_2
  CLASS  CORE ;
  FOREIGN sdffnh_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 28.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 24.000 8.450 26.000 9.050 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 16.950 0.000 17.550 2.700 ;
        RECT 0.000 0.000 28.750 2.500 ;
    END
  END vss!
  PIN ckb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 26.500 8.450 28.500 9.050 ;
    END
  END ckb
  PIN se
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.100 8.350 8.650 9.150 ;
    END
  END se
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.450 8.350 3.000 9.150 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 3.450 13.550 4.050 16.250 ;
        RECT 0.000 13.750 28.750 16.250 ;
        RECT 23.350 13.500 23.950 16.250 ;
        RECT 17.250 13.550 17.850 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 21.500 8.450 23.500 9.050 ;
    END
  END qb
  PIN g
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.850 6.450 3.450 7.800 ;
        RECT 3.500 8.450 5.300 9.050 ;
        RECT 3.500 7.200 4.100 9.050 ;
        RECT 2.850 7.200 4.100 7.800 ;
    END
  END g
  PIN sdi
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 10.250 8.350 12.000 9.100 ;
    END
  END sdi
  OBS 
      LAYER Metal1 ;
        RECT 6.000 5.900 8.600 6.500 ;
        RECT 0.350 6.050 0.950 10.300 ;
        RECT 6.000 5.900 6.600 10.300 ;
        RECT 0.350 9.700 6.750 10.300 ;
        RECT 9.700 6.900 10.300 7.800 ;
        RECT 9.150 7.200 12.000 7.800 ;
        RECT 9.150 7.200 9.750 10.300 ;
        RECT 8.250 9.700 9.750 10.300 ;
        RECT 12.500 5.900 14.250 6.500 ;
        RECT 12.500 5.900 13.100 10.300 ;
        RECT 12.500 9.700 15.450 10.300 ;
        RECT 15.550 6.600 19.600 7.200 ;
        RECT 15.550 6.600 16.250 7.950 ;
        RECT 13.600 7.300 16.250 7.950 ;
        RECT 4.900 4.800 23.350 5.400 ;
        RECT 22.750 4.800 23.350 6.750 ;
        RECT 4.900 4.800 5.500 7.600 ;
        RECT 20.300 7.250 28.400 7.850 ;
        RECT 17.550 7.700 18.150 9.200 ;
        RECT 20.300 7.250 20.900 9.200 ;
        RECT 13.850 8.600 20.900 9.200 ;
  END 
END sdffnh_2

MACRO sdffnh_1
  CLASS  CORE ;
  FOREIGN sdffnh_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 28.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 26.500 5.950 28.500 6.550 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 3.350 0.000 3.950 2.700 ;
        RECT 0.000 0.000 28.750 2.500 ;
        RECT 25.400 0.000 26.000 2.700 ;
        RECT 6.200 0.000 6.800 2.700 ;
    END
  END vss!
  PIN ckb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 15.450 3.450 18.900 4.050 ;
    END
  END ckb
  PIN se
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.750 8.450 7.750 9.050 ;
    END
  END se
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.450 8.400 3.300 9.100 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 3.450 13.550 4.050 16.250 ;
        RECT 0.000 13.750 28.750 16.250 ;
        RECT 25.400 13.550 26.000 16.250 ;
        RECT 17.400 13.550 18.000 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 24.700 8.450 26.700 9.050 ;
    END
  END qb
  PIN g
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.350 5.950 4.050 7.800 ;
        RECT 3.800 7.200 4.400 9.050 ;
    END
  END g
  PIN sdi
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 10.200 8.450 12.250 9.050 ;
    END
  END sdi
  OBS 
      LAYER Metal1 ;
        RECT 0.350 5.950 0.950 10.300 ;
        RECT 0.350 9.700 6.750 10.300 ;
        RECT 0.350 3.450 6.750 4.050 ;
        RECT 6.150 5.950 8.600 6.550 ;
        RECT 9.700 6.900 10.300 7.800 ;
        RECT 9.100 7.200 12.200 7.800 ;
        RECT 9.100 7.200 9.700 9.200 ;
        RECT 8.250 8.600 9.700 9.200 ;
        RECT 12.750 5.950 14.400 6.550 ;
        RECT 12.750 5.950 13.350 10.250 ;
        RECT 12.750 9.650 15.000 10.250 ;
        RECT 14.750 8.350 15.350 9.050 ;
        RECT 14.750 8.450 22.250 9.050 ;
        RECT 13.850 7.050 14.450 7.850 ;
        RECT 21.200 7.150 22.250 7.750 ;
        RECT 13.850 7.250 16.750 7.850 ;
        RECT 15.850 7.350 21.800 7.950 ;
        RECT 22.400 6.000 23.500 6.600 ;
        RECT 22.900 6.000 23.500 10.300 ;
        RECT 21.900 9.700 23.500 10.300 ;
  END 
END sdffnh_1

MACRO sdffn_8
  CLASS  CORE ;
  FOREIGN sdffn_8 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 31.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 25.950 8.450 27.950 9.050 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 3.400 0.000 4.000 2.650 ;
        RECT 0.000 0.000 31.250 2.500 ;
    END
  END vss!
  PIN ckb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 28.700 4.700 30.700 5.300 ;
    END
  END ckb
  PIN se
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.450 5.800 4.050 9.050 ;
        RECT 3.450 5.800 5.150 6.400 ;
        RECT 2.100 8.400 4.050 9.050 ;
    END
  END se
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.800 5.950 2.800 6.550 ;
        RECT 2.200 5.950 2.800 6.950 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 3.400 13.450 4.000 16.250 ;
        RECT 0.000 13.750 31.250 16.250 ;
        RECT 21.500 13.450 22.100 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 21.800 8.450 24.050 9.050 ;
    END
  END qb
  PIN sdi
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.250 8.450 5.850 10.300 ;
        RECT 4.700 9.700 5.850 10.300 ;
    END
  END sdi
  OBS 
      LAYER Metal1 ;
        RECT 0.450 4.700 6.950 5.300 ;
        RECT 6.350 4.700 6.950 10.100 ;
        RECT 7.900 5.150 9.150 5.750 ;
        RECT 7.900 5.150 8.500 10.300 ;
        RECT 7.900 9.700 9.150 10.300 ;
        RECT 11.200 7.200 17.150 7.800 ;
        RECT 16.550 7.200 17.150 7.850 ;
        RECT 11.200 7.200 11.800 8.500 ;
        RECT 10.500 7.900 11.800 8.500 ;
        RECT 18.500 7.050 19.100 9.050 ;
        RECT 15.400 8.450 19.100 9.050 ;
        RECT 13.450 9.000 14.050 10.300 ;
        RECT 13.450 9.700 20.400 10.300 ;
        RECT 15.150 4.700 25.900 5.300 ;
        RECT 9.650 5.950 22.350 6.550 ;
        RECT 9.000 6.350 10.250 6.950 ;
        RECT 21.750 5.950 22.350 7.800 ;
        RECT 21.750 7.200 30.600 7.800 ;
        RECT 9.000 6.350 9.600 9.000 ;
  END 
END sdffn_8

MACRO sdffn_6
  CLASS  CORE ;
  FOREIGN sdffn_6 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 30.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 24.600 9.700 26.600 10.300 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 3.050 0.000 3.650 2.800 ;
        RECT 0.000 0.000 30.000 2.500 ;
        RECT 23.800 0.000 24.400 2.650 ;
    END
  END vss!
  PIN ckb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 27.500 5.950 29.500 6.550 ;
    END
  END ckb
  PIN se
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.450 6.450 4.050 9.050 ;
        RECT 3.450 6.450 4.600 7.100 ;
        RECT 2.200 8.450 4.050 9.050 ;
    END
  END se
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.400 5.950 2.400 6.550 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 3.400 13.450 4.000 16.250 ;
        RECT 0.000 13.750 30.000 16.250 ;
        RECT 23.800 13.450 24.400 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 19.100 8.450 21.100 9.050 ;
    END
  END qb
  PIN sdi
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.500 4.700 5.500 5.300 ;
    END
  END sdi
  OBS 
      LAYER Metal1 ;
        RECT 0.450 9.700 6.950 10.300 ;
        RECT 7.600 4.850 8.800 5.450 ;
        RECT 7.600 4.850 8.200 10.400 ;
        RECT 7.600 9.800 8.800 10.400 ;
        RECT 13.200 6.050 13.800 7.800 ;
        RECT 10.050 7.200 13.800 7.800 ;
        RECT 11.950 9.650 22.700 10.250 ;
        RECT 14.300 5.900 15.050 6.500 ;
        RECT 14.450 7.100 24.000 7.700 ;
        RECT 14.450 5.900 15.050 8.900 ;
        RECT 9.950 4.700 25.750 5.300 ;
        RECT 15.600 4.700 16.200 5.750 ;
        RECT 9.950 4.700 10.550 6.550 ;
        RECT 8.700 5.950 10.550 6.550 ;
        RECT 25.150 4.700 25.750 7.800 ;
        RECT 25.150 7.200 29.550 7.800 ;
        RECT 8.700 5.950 9.300 8.900 ;
        RECT 8.700 8.300 13.750 8.900 ;
  END 
END sdffn_6

MACRO sdffn_4
  CLASS  CORE ;
  FOREIGN sdffn_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 30.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 25.550 7.200 27.550 7.800 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 30.000 2.500 ;
    END
  END vss!
  PIN ckb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 12.450 5.950 14.450 6.550 ;
    END
  END ckb
  PIN se
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.350 5.650 1.550 6.250 ;
        RECT 0.950 8.400 2.200 9.000 ;
        RECT 0.950 5.650 1.550 9.000 ;
    END
  END se
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.000 6.450 3.600 7.800 ;
        RECT 3.000 7.200 4.700 7.800 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 30.000 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 21.250 5.950 23.250 6.550 ;
    END
  END qb
  PIN sdi
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.350 8.450 7.350 9.050 ;
    END
  END sdi
  OBS 
      LAYER Metal1 ;
        RECT 5.200 6.200 8.050 6.800 ;
        RECT 9.000 6.200 10.050 6.800 ;
        RECT 9.000 6.200 9.600 7.950 ;
        RECT 8.250 7.350 9.600 7.950 ;
        RECT 8.250 7.350 8.850 10.250 ;
        RECT 8.250 9.650 10.050 10.250 ;
        RECT 19.400 6.800 20.000 7.950 ;
        RECT 10.250 7.350 20.000 7.950 ;
        RECT 9.350 8.450 20.450 9.050 ;
  END 
END sdffn_4

MACRO sdffn_3
  CLASS  CORE ;
  FOREIGN sdffn_3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 27.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 23.550 5.950 25.550 6.550 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 27.500 2.500 ;
    END
  END vss!
  PIN ckb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 12.950 5.950 14.950 6.550 ;
    END
  END ckb
  PIN se
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.350 6.250 0.950 7.300 ;
        RECT 0.350 6.700 2.800 7.300 ;
        RECT 0.350 6.550 1.650 7.300 ;
        RECT 0.950 6.550 1.550 7.800 ;
    END
  END se
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.450 6.800 4.100 9.050 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 27.500 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 20.250 5.950 22.250 6.550 ;
    END
  END qb
  PIN sdi
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.950 8.000 6.550 10.400 ;
    END
  END sdi
  OBS 
      LAYER Metal1 ;
        RECT 5.150 6.250 8.000 6.850 ;
        RECT 9.100 6.050 10.050 6.650 ;
        RECT 9.100 6.050 9.700 7.950 ;
        RECT 8.200 7.350 9.700 7.950 ;
        RECT 8.200 7.350 8.800 10.150 ;
        RECT 8.200 9.550 10.050 10.150 ;
        RECT 9.300 8.450 19.600 9.050 ;
        RECT 10.200 7.350 19.650 7.950 ;
  END 
END sdffn_3

MACRO sdffn_2
  CLASS  CORE ;
  FOREIGN sdffn_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 23.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 19.000 8.450 21.000 9.050 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 11.600 0.000 12.200 2.700 ;
        RECT 0.000 0.000 23.750 2.500 ;
        RECT 17.600 0.000 18.200 2.800 ;
    END
  END vss!
  PIN ckb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 21.500 8.450 23.500 9.050 ;
    END
  END ckb
  PIN se
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.450 6.450 4.050 7.100 ;
        RECT 3.450 5.950 4.050 9.050 ;
    END
  END se
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.700 6.250 5.300 8.750 ;
        RECT 4.700 7.200 5.550 7.800 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 11.900 13.550 12.500 16.250 ;
        RECT 0.000 13.750 23.750 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 16.150 8.450 18.150 9.050 ;
    END
  END qb
  PIN sdi
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.350 8.350 2.950 9.100 ;
    END
  END sdi
  OBS 
      LAYER Metal1 ;
        RECT 0.250 6.300 0.850 10.300 ;
        RECT 6.050 5.850 6.650 10.300 ;
        RECT 0.250 9.700 6.650 10.300 ;
        RECT 7.150 5.850 8.850 6.450 ;
        RECT 7.150 5.850 7.750 10.150 ;
        RECT 7.150 9.550 9.200 10.150 ;
        RECT 8.400 7.050 9.000 7.950 ;
        RECT 10.250 6.900 14.200 7.500 ;
        RECT 8.400 7.350 10.900 7.950 ;
        RECT 14.750 7.250 23.400 7.850 ;
        RECT 12.200 8.000 15.350 8.600 ;
        RECT 14.750 7.250 15.350 8.600 ;
        RECT 8.250 8.450 12.800 9.050 ;
  END 
END sdffn_2

MACRO or3i_5
  CLASS  CORE ;
  FOREIGN or3i_5 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.000 5.950 5.000 6.550 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 13.750 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.000 5.950 10.000 6.550 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 11.200 9.700 13.200 10.300 ;
    END
  END c
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 3.350 13.600 3.950 16.250 ;
        RECT 0.000 13.750 13.750 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.150 9.700 6.150 10.300 ;
    END
  END x
END or3i_5

MACRO or3i_4
  CLASS  CORE ;
  FOREIGN or3i_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.600 5.950 2.600 6.550 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 11.250 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.250 7.200 10.250 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.500 5.950 10.500 6.550 ;
    END
  END c
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 11.250 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.350 7.200 4.050 7.800 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 4.500 5.900 8.000 6.600 ;
  END 
END or3i_4

MACRO or3i_3
  CLASS  CORE ;
  FOREIGN or3i_3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.900 5.950 4.900 6.550 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 10.000 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.900 5.950 7.900 6.550 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.250 8.450 9.250 9.050 ;
    END
  END c
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 4.100 13.550 4.850 16.250 ;
        RECT 0.000 13.750 10.000 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.750 8.450 3.750 9.050 ;
    END
  END x
END or3i_3

MACRO or3i_2
  CLASS  CORE ;
  FOREIGN or3i_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.900 5.950 2.900 6.550 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 7.500 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.950 7.200 4.950 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.100 8.450 7.100 9.050 ;
    END
  END c
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 7.500 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.350 8.450 2.750 9.050 ;
    END
  END x
END or3i_2

MACRO or3i_1
  CLASS  CORE ;
  FOREIGN or3i_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.900 5.950 2.900 6.550 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 7.500 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.350 7.200 5.350 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.100 8.450 7.100 9.050 ;
    END
  END c
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 7.500 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.350 8.450 2.750 9.050 ;
    END
  END x
END or3i_1

MACRO or3_5
  CLASS  CORE ;
  FOREIGN or3_5 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.150 5.950 10.150 6.550 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 3.050 0.000 3.650 2.550 ;
        RECT 0.000 0.000 12.500 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.700 5.650 6.300 6.550 ;
        RECT 5.700 5.950 7.650 6.550 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.950 5.950 4.950 6.650 ;
    END
  END c
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 12.500 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.450 5.950 2.450 6.550 ;
    END
  END x
END or3_5

MACRO or3_4
  CLASS  CORE ;
  FOREIGN or3_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.750 7.200 9.750 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 7.300 0.000 8.000 2.700 ;
        RECT 0.000 0.000 10.000 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.550 5.950 7.550 6.550 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.700 5.950 4.700 6.550 ;
    END
  END c
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.450 13.650 1.050 16.250 ;
        RECT 0.000 13.750 10.000 16.250 ;
        RECT 3.550 13.500 4.250 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.500 7.200 2.500 7.800 ;
    END
  END x
END or3_4

MACRO or3_3
  CLASS  CORE ;
  FOREIGN or3_3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.600 8.450 9.600 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 10.000 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.950 7.050 6.550 9.050 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.100 8.450 5.100 9.050 ;
    END
  END c
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 10.000 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.400 5.950 3.400 6.550 ;
    END
  END x
END or3_3

MACRO or3_2
  CLASS  CORE ;
  FOREIGN or3_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.100 8.450 7.100 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 7.500 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.350 7.200 5.350 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.900 8.450 2.900 9.050 ;
    END
  END c
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 2.100 13.550 2.800 16.250 ;
        RECT 0.000 13.750 7.500 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.400 5.950 2.400 6.550 ;
    END
  END x
END or3_2

MACRO or3_1
  CLASS  CORE ;
  FOREIGN or3_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.100 8.450 7.100 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 7.500 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.450 7.200 5.450 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.400 8.450 3.400 9.050 ;
    END
  END c
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 7.500 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.350 5.950 2.350 6.550 ;
    END
  END x
END or3_1

MACRO or2_8
  CLASS  CORE ;
  FOREIGN or2_8 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.900 7.200 2.900 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 12.500 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.500 8.450 2.500 9.100 ;
        RECT 1.500 8.450 6.600 9.050 ;
        RECT 5.300 8.400 5.900 9.050 ;
    END
  END b
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 9.350 13.550 10.050 16.250 ;
        RECT 0.000 13.750 12.500 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.650 8.450 11.700 9.050 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 3.400 7.200 10.700 7.800 ;
  END 
END or2_8

MACRO or2_6
  CLASS  CORE ;
  FOREIGN or2_6 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.550 7.200 2.550 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 4.750 0.000 5.350 2.600 ;
        RECT 0.000 0.000 10.000 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.200 8.450 2.500 9.100 ;
        RECT 1.200 8.450 5.400 9.050 ;
    END
  END b
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 10.000 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.150 8.450 9.150 9.050 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 3.050 7.200 8.950 7.800 ;
  END 
END or2_6

MACRO or2_5
  CLASS  CORE ;
  FOREIGN or2_5 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.550 7.200 2.550 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 10.000 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.150 8.450 2.200 9.100 ;
        RECT 1.150 8.450 5.350 9.050 ;
    END
  END b
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 10.000 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.150 8.450 9.150 9.050 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 3.050 7.200 8.950 7.800 ;
  END 
END or2_5

MACRO or2_4
  CLASS  CORE ;
  FOREIGN or2_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.550 7.000 2.150 9.050 ;
        RECT 0.950 8.450 2.150 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 7.500 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.900 8.150 3.500 9.050 ;
        RECT 2.650 8.350 4.250 9.050 ;
    END
  END b
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 7.500 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.750 8.450 5.350 10.450 ;
        RECT 4.750 8.450 7.050 9.050 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 0.450 5.800 4.650 6.400 ;
        RECT 4.050 5.800 4.650 7.600 ;
        RECT 0.450 5.800 1.050 7.600 ;
        RECT 4.050 7.000 5.200 7.600 ;
  END 
END or2_4

MACRO or2_3
  CLASS  CORE ;
  FOREIGN or2_3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 8.400 2.050 9.100 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 7.500 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.550 8.350 4.250 9.100 ;
    END
  END b
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 3.050 13.550 3.650 16.250 ;
        RECT 0.000 13.750 7.500 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.750 8.400 7.000 9.100 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 2.150 6.250 2.750 7.800 ;
        RECT 2.150 7.200 5.050 7.800 ;
  END 
END or2_3

MACRO or2_2
  CLASS  CORE ;
  FOREIGN or2_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 8.400 2.050 9.100 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 6.250 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.550 8.400 4.350 9.100 ;
    END
  END b
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 3.050 13.550 3.750 16.250 ;
        RECT 0.000 13.750 6.250 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.700 5.950 5.450 6.550 ;
        RECT 4.850 5.950 5.450 9.100 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 1.250 7.200 4.100 7.800 ;
  END 
END or2_2

MACRO or2_1
  CLASS  CORE ;
  FOREIGN or2_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 8.400 2.000 9.100 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 6.250 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.500 8.450 4.500 9.050 ;
    END
  END b
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 3.100 13.550 3.700 16.250 ;
        RECT 0.000 13.750 6.250 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.800 5.950 5.800 6.550 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 1.350 7.200 4.250 7.800 ;
  END 
END or2_1

MACRO oaoi211_5
  CLASS  CORE ;
  FOREIGN oaoi211_5 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 25.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 13.450 5.950 24.050 6.550 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 19.650 0.000 20.250 2.700 ;
        RECT 0.000 0.000 25.000 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 11.650 7.050 12.600 7.850 ;
        RECT 11.650 7.250 22.700 7.850 ;
        RECT 11.650 7.200 15.300 7.850 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.150 7.100 10.550 7.800 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.350 4.700 5.350 5.300 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 25.000 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.750 5.950 9.850 6.550 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 7.550 3.450 21.950 4.050 ;
        RECT 2.450 9.700 24.550 10.300 ;
  END 
END oaoi211_5

MACRO oaoi211_4
  CLASS  CORE ;
  FOREIGN oaoi211_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 22.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 12.050 5.950 20.400 6.550 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 22.500 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 11.500 7.200 21.100 7.850 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.900 7.200 10.350 7.800 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.850 7.200 5.750 7.850 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 22.500 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.650 5.950 9.750 6.550 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 2.350 9.700 19.250 10.300 ;
        RECT 7.450 3.450 21.850 4.050 ;
  END 
END oaoi211_4

MACRO oaoi211_3
  CLASS  CORE ;
  FOREIGN oaoi211_3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 22.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 12.050 7.150 15.300 7.750 ;
        RECT 14.700 7.200 20.300 7.800 ;
        RECT 18.750 7.150 20.300 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 22.500 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 11.500 8.450 21.100 9.050 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.750 8.450 10.450 9.050 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.750 8.450 5.750 9.050 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 22.500 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.650 7.200 9.750 7.800 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 7.450 4.700 18.350 5.300 ;
        RECT 2.350 9.700 19.250 10.300 ;
  END 
END oaoi211_3

MACRO oaoi211_2
  CLASS  CORE ;
  FOREIGN oaoi211_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 16.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.850 8.450 13.800 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 16.250 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.700 7.200 15.300 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.650 8.450 6.650 9.050 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 8.450 2.250 9.050 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 16.250 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.300 7.200 5.450 7.800 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 0.450 9.700 13.050 10.300 ;
        RECT 3.850 4.700 14.750 5.300 ;
  END 
END oaoi211_2

MACRO oaoi211_1
  CLASS  CORE ;
  FOREIGN oaoi211_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.300 7.200 12.300 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 13.750 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 10.500 8.450 12.800 9.050 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.650 8.450 6.650 9.050 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.850 8.450 3.900 9.050 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 13.750 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.150 5.950 6.150 6.550 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 7.250 5.950 11.250 6.550 ;
        RECT 0.450 9.700 13.050 10.300 ;
  END 
END oaoi211_1

MACRO oai33_6
  CLASS  CORE ;
  FOREIGN oai33_6 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 33.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 14.700 8.150 15.300 9.050 ;
        RECT 1.200 8.400 15.300 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 3.750 0.000 4.350 2.800 ;
        RECT 0.000 0.000 33.750 2.500 ;
        RECT 13.900 0.000 14.600 2.750 ;
        RECT 7.100 0.000 7.800 2.750 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.400 5.950 1.250 6.700 ;
        RECT 0.400 5.950 9.900 6.550 ;
        RECT 6.250 5.950 7.300 6.700 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.700 7.200 14.050 7.800 ;
        RECT 17.200 7.050 17.800 8.250 ;
        RECT 13.450 7.050 17.800 7.650 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 24.850 5.950 28.300 6.550 ;
        RECT 27.700 5.950 28.300 8.250 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 29.050 7.200 31.050 7.850 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 33.750 16.250 ;
    END
  END vdd!
  PIN f
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 18.700 7.100 23.150 7.700 ;
        RECT 25.950 8.750 31.800 9.350 ;
        RECT 31.200 8.400 31.800 9.350 ;
        RECT 22.550 8.450 26.550 9.050 ;
        RECT 25.300 8.200 26.550 9.050 ;
        RECT 22.550 8.350 23.550 9.050 ;
        RECT 22.550 7.100 23.150 9.050 ;
    END
  END f
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 21.400 8.450 22.050 10.300 ;
        RECT 23.750 9.850 29.050 10.450 ;
        RECT 0.450 9.700 24.850 10.300 ;
        RECT 21.400 9.600 22.150 10.300 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 19.200 5.800 24.300 6.400 ;
        RECT 23.700 5.800 24.300 7.800 ;
        RECT 2.050 3.450 29.850 4.050 ;
  END 
END oai33_6

MACRO oai33_5
  CLASS  CORE ;
  FOREIGN oai33_5 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 27.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.550 7.300 7.550 9.350 ;
        RECT 6.550 8.750 15.100 9.350 ;
        RECT 14.500 6.200 15.100 9.350 ;
        RECT 11.900 6.200 15.100 6.800 ;
        RECT 0.300 8.500 7.800 9.100 ;
        RECT 6.550 8.450 7.800 9.350 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 4.800 0.000 5.500 2.700 ;
        RECT 0.000 0.000 27.500 2.500 ;
        RECT 11.650 0.000 12.250 2.800 ;
        RECT 8.250 0.000 8.850 2.800 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.450 7.200 3.450 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.950 5.950 4.600 8.000 ;
        RECT 10.550 5.950 11.150 7.150 ;
        RECT 10.300 5.950 11.150 6.650 ;
        RECT 1.250 5.950 11.150 6.550 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 15.950 7.100 16.550 9.050 ;
        RECT 15.950 8.450 24.300 9.050 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 18.000 6.350 18.600 7.800 ;
        RECT 18.000 7.200 25.550 7.800 ;
        RECT 20.000 7.100 21.600 7.800 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 27.500 16.250 ;
    END
  END vdd!
  PIN f
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 19.250 5.950 27.050 6.550 ;
    END
  END f
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.450 9.850 17.800 10.450 ;
        RECT 17.200 9.700 23.000 10.300 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 9.250 7.250 9.950 8.250 ;
        RECT 13.200 7.300 13.800 8.250 ;
        RECT 9.250 7.650 13.800 8.250 ;
        RECT 3.150 3.450 24.500 4.050 ;
  END 
END oai33_5

MACRO oai33_4
  CLASS  CORE ;
  FOREIGN oai33_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 23.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 11.450 6.700 12.050 9.050 ;
        RECT 4.250 8.450 12.050 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 23.750 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.450 5.950 4.050 6.850 ;
        RECT 7.450 5.950 8.050 6.750 ;
        RECT 3.450 5.950 8.050 6.550 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.950 7.200 1.550 8.000 ;
        RECT 0.950 7.350 10.050 7.950 ;
        RECT 9.450 6.700 10.050 7.950 ;
        RECT 0.950 7.350 2.300 8.000 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 14.850 7.050 15.450 9.050 ;
        RECT 14.850 8.450 20.550 9.050 ;
        RECT 14.850 8.300 15.950 9.050 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 18.000 7.150 19.050 7.900 ;
        RECT 18.000 7.300 22.300 7.900 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 15.700 13.450 16.300 16.250 ;
        RECT 0.000 13.750 23.750 16.250 ;
    END
  END vdd!
  PIN f
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 16.450 5.950 17.100 7.650 ;
        RECT 16.450 5.950 23.400 6.550 ;
    END
  END f
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 13.450 5.850 14.050 10.300 ;
        RECT 5.200 9.700 19.800 10.300 ;
        RECT 13.450 5.850 14.550 6.450 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 2.050 3.450 23.050 4.050 ;
  END 
END oai33_4

MACRO oai33_3
  CLASS  CORE ;
  FOREIGN oai33_3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 20.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.200 8.450 7.400 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.350 0.000 0.950 2.800 ;
        RECT 0.000 0.000 20.000 2.500 ;
        RECT 7.200 0.000 7.800 2.800 ;
        RECT 3.800 0.000 4.400 2.800 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.700 7.200 8.400 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.050 5.800 2.650 7.950 ;
        RECT 8.900 7.100 11.200 7.800 ;
        RECT 10.600 6.800 11.200 7.800 ;
        RECT 8.900 5.800 9.500 7.800 ;
        RECT 2.050 5.800 9.500 6.400 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 15.300 7.200 16.200 8.200 ;
        RECT 14.700 7.200 18.450 7.800 ;
        RECT 17.850 7.150 18.450 7.800 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 10.000 5.700 14.150 6.300 ;
        RECT 13.350 6.000 15.050 6.600 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 4.050 13.450 4.650 16.250 ;
        RECT 0.000 13.750 20.000 16.250 ;
    END
  END vdd!
  PIN f
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 12.100 7.000 12.700 9.300 ;
        RECT 17.100 8.450 18.200 9.050 ;
        RECT 12.100 8.700 17.900 9.300 ;
    END
  END f
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.450 9.700 9.050 10.300 ;
        RECT 8.450 9.800 19.650 10.400 ;
        RECT 19.050 5.700 19.650 10.400 ;
        RECT 15.550 5.700 19.650 6.300 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 2.050 4.600 17.850 5.200 ;
  END 
END oai33_3

MACRO oai33_2
  CLASS  CORE ;
  FOREIGN oai33_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 16.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.450 7.200 3.800 7.800 ;
        RECT 2.850 7.200 3.800 7.850 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.950 0.000 1.550 2.800 ;
        RECT 0.000 0.000 16.250 2.500 ;
        RECT 8.400 0.000 9.000 2.950 ;
        RECT 5.000 0.000 5.600 2.950 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.300 5.950 6.000 6.550 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.650 5.850 7.300 9.050 ;
        RECT 1.200 8.450 7.300 9.050 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.850 5.950 10.450 7.600 ;
        RECT 9.850 5.950 15.800 6.550 ;
        RECT 9.850 5.950 10.950 6.650 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 11.400 7.200 13.700 7.800 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 16.250 16.250 ;
    END
  END vdd!
  PIN f
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.800 7.350 8.400 9.050 ;
        RECT 13.450 8.450 14.300 9.100 ;
        RECT 7.800 8.450 14.300 9.050 ;
    END
  END f
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.950 9.700 11.600 10.300 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 3.300 3.450 14.100 4.050 ;
  END 
END oai33_2

MACRO oai33_1
  CLASS  CORE ;
  FOREIGN oai33_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.350 7.200 3.700 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 12.500 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.200 7.200 6.200 7.900 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.200 8.450 7.250 9.050 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.650 5.950 11.650 6.550 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.850 7.200 10.850 7.800 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 12.500 16.250 ;
    END
  END vdd!
  PIN f
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.550 6.200 8.350 6.800 ;
        RECT 7.750 8.450 9.150 9.100 ;
        RECT 7.750 6.200 8.350 9.100 ;
        RECT 7.100 6.200 8.350 7.200 ;
    END
  END f
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.950 9.700 12.050 10.300 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 2.100 3.450 9.950 4.050 ;
  END 
END oai33_1

MACRO oai31_6
  CLASS  CORE ;
  FOREIGN oai31_6 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 22.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.650 7.750 5.250 9.050 ;
        RECT 4.650 8.450 20.300 9.050 ;
        RECT 10.300 7.400 10.900 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 11.900 0.000 12.600 2.750 ;
        RECT 0.000 0.000 22.500 2.500 ;
        RECT 15.350 0.000 15.950 2.800 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 12.700 7.200 17.800 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 14.600 5.950 16.600 6.550 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.350 7.200 2.350 7.800 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 7.300 13.550 8.000 16.250 ;
        RECT 0.000 13.750 22.500 16.250 ;
        RECT 14.300 13.550 15.000 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.900 6.250 3.500 10.300 ;
        RECT 0.450 9.700 18.450 10.300 ;
        RECT 2.900 6.250 4.450 7.200 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 2.150 4.700 21.050 5.300 ;
  END 
END oai31_6

MACRO oai31_5
  CLASS  CORE ;
  FOREIGN oai31_5 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 20.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.950 7.200 5.550 9.050 ;
        RECT 4.950 8.450 18.050 9.050 ;
        RECT 10.300 8.350 11.050 9.050 ;
        RECT 10.450 7.400 11.050 9.050 ;
        RECT 4.950 8.350 6.050 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 15.350 0.000 15.950 2.800 ;
        RECT 0.000 0.000 20.000 2.500 ;
        RECT 18.750 0.000 19.350 2.800 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 13.050 6.750 13.650 7.800 ;
        RECT 13.050 7.200 19.050 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 14.600 5.950 16.600 6.550 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.350 7.200 3.350 7.800 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 7.650 13.550 8.350 16.250 ;
        RECT 0.000 13.750 20.000 16.250 ;
        RECT 14.650 13.550 15.350 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.850 5.850 4.450 10.300 ;
        RECT 0.450 9.700 18.800 10.300 ;
        RECT 3.850 9.600 4.600 10.300 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 2.150 4.700 17.650 5.300 ;
  END 
END oai31_5

MACRO oai31_4
  CLASS  CORE ;
  FOREIGN oai31_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 18.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.250 8.450 17.550 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 5.700 0.000 6.300 2.800 ;
        RECT 0.000 0.000 18.750 2.500 ;
        RECT 12.500 0.000 13.100 2.800 ;
        RECT 9.100 0.000 9.700 2.800 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.450 7.200 16.450 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 12.500 5.950 14.500 6.550 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.800 8.450 2.800 9.050 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 7.150 13.550 7.850 16.250 ;
        RECT 0.000 13.750 18.750 16.250 ;
        RECT 14.150 13.550 14.850 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.450 9.700 18.300 10.300 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 3.700 4.700 14.800 5.300 ;
  END 
END oai31_4

MACRO oai31_3
  CLASS  CORE ;
  FOREIGN oai31_3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.850 6.550 4.450 9.050 ;
        RECT 3.850 8.450 11.000 9.050 ;
        RECT 10.300 8.300 11.000 9.050 ;
        RECT 3.850 8.350 4.600 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 6.700 0.000 7.400 2.700 ;
        RECT 0.000 0.000 15.000 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.250 5.950 8.850 6.600 ;
        RECT 8.250 5.950 10.250 6.550 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 12.500 7.200 14.500 7.800 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.600 7.200 2.600 7.800 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 6.550 13.550 7.250 16.250 ;
        RECT 0.000 13.750 15.000 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.200 9.700 10.700 10.300 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 0.350 4.700 12.450 5.300 ;
  END 
END oai31_3

MACRO oai31_2
  CLASS  CORE ;
  FOREIGN oai31_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.800 5.950 6.800 6.550 ;
        RECT 6.200 5.950 6.800 6.650 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 3.850 0.000 4.450 2.800 ;
        RECT 0.000 0.000 11.250 2.500 ;
        RECT 10.300 0.000 10.900 2.750 ;
        RECT 7.350 0.000 7.950 2.650 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.300 7.200 9.050 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.950 7.550 3.550 9.050 ;
        RECT 2.950 8.450 10.300 9.050 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.450 7.200 2.450 7.800 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 11.250 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.450 9.700 6.750 10.300 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 2.150 4.700 9.550 5.300 ;
  END 
END oai31_2

MACRO oai31_1
  CLASS  CORE ;
  FOREIGN oai31_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.400 7.200 7.400 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 11.250 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.900 7.200 9.900 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.050 7.200 4.050 7.800 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.950 5.950 2.950 6.550 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 11.250 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.750 8.450 6.650 9.050 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 2.550 4.700 7.550 5.300 ;
  END 
END oai31_1

MACRO oai22_6
  CLASS  CORE ;
  FOREIGN oai22_6 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 22.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 12.900 7.200 14.850 7.850 ;
        RECT 12.900 7.200 21.550 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 22.500 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 11.800 5.950 21.500 6.550 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.100 7.200 5.400 7.800 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.700 7.200 10.700 7.800 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 5.650 13.550 6.350 16.250 ;
        RECT 0.000 13.750 22.500 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.100 9.700 19.350 10.300 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 0.500 4.700 21.500 5.300 ;
  END 
END oai22_6

MACRO oai22_5
  CLASS  CORE ;
  FOREIGN oai22_5 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 20.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 11.450 7.200 17.500 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 20.000 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.300 5.950 19.550 6.550 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 5.800 1.900 6.550 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.350 7.200 8.350 7.800 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 3.150 13.550 3.850 16.250 ;
        RECT 0.000 13.750 20.000 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.600 9.700 16.850 10.300 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 2.400 5.850 6.400 6.450 ;
        RECT 0.700 4.700 18.450 5.300 ;
  END 
END oai22_5

MACRO oai22_4
  CLASS  CORE ;
  FOREIGN oai22_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 17.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 11.450 7.200 16.550 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 9.200 0.000 9.800 2.700 ;
        RECT 0.000 0.000 17.500 2.500 ;
        RECT 12.700 0.000 13.300 2.700 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.650 5.950 13.350 6.550 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.850 7.200 2.850 7.800 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.850 7.200 7.850 7.800 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 3.150 13.550 3.850 16.250 ;
        RECT 0.000 13.750 17.500 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.600 9.700 16.850 10.300 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 0.700 4.700 15.050 5.300 ;
  END 
END oai22_4

MACRO oai22_3
  CLASS  CORE ;
  FOREIGN oai22_3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.250 8.450 14.050 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 15.000 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.650 7.200 11.650 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.800 7.200 2.800 7.850 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.150 5.950 7.150 6.550 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 15.000 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.300 9.700 14.350 10.300 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 0.350 4.700 11.200 5.300 ;
  END 
END oai22_3

MACRO oai22_2
  CLASS  CORE ;
  FOREIGN oai22_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.800 8.450 10.500 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 12.500 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.350 7.200 7.200 7.850 ;
        RECT 6.350 7.200 11.000 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.400 7.150 5.350 7.850 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.450 7.200 2.800 7.800 ;
        RECT 1.550 7.200 2.800 7.850 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 12.500 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.300 9.700 9.150 10.300 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 1.650 4.700 9.350 5.300 ;
  END 
END oai22_2

MACRO oai22_1
  CLASS  CORE ;
  FOREIGN oai22_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.750 7.200 7.800 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 8.750 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.000 8.450 7.600 10.300 ;
        RECT 7.000 9.700 8.050 10.300 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 7.200 1.600 7.800 ;
        RECT 1.000 7.200 1.600 8.700 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.250 7.200 5.250 7.800 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 8.750 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.150 7.150 2.750 10.300 ;
        RECT 0.400 9.700 5.700 10.300 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 0.450 4.700 7.850 5.300 ;
  END 
END oai22_1

MACRO oai222_5
  CLASS  CORE ;
  FOREIGN oai222_5 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 31.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 14.650 8.450 19.650 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 9.550 0.000 10.250 2.750 ;
        RECT 0.000 0.000 31.250 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 12.100 7.200 12.800 9.100 ;
        RECT 12.100 7.200 16.550 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 23.300 7.000 29.600 7.600 ;
        RECT 28.450 7.200 30.400 7.800 ;
        RECT 28.950 7.000 29.600 8.900 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 22.550 8.100 23.350 9.050 ;
        RECT 22.100 8.450 27.100 9.050 ;
        RECT 26.450 8.100 27.100 9.050 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.250 8.450 9.250 9.050 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 31.250 16.250 ;
    END
  END vdd!
  PIN f
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.700 7.200 2.300 9.100 ;
        RECT 1.700 7.200 7.700 7.800 ;
    END
  END f
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 21.000 5.800 21.600 10.300 ;
        RECT 3.600 9.700 30.350 10.300 ;
        RECT 21.000 5.800 28.450 6.400 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 6.100 5.800 10.200 6.400 ;
        RECT 4.400 4.700 18.700 5.300 ;
        RECT 19.750 4.700 30.150 5.300 ;
        RECT 19.750 4.700 20.350 6.400 ;
        RECT 12.900 5.800 20.350 6.400 ;
  END 
END oai222_5

MACRO oai222_4
  CLASS  CORE ;
  FOREIGN oai222_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 25.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.100 7.200 13.450 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 25.000 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 10.850 8.450 16.000 9.050 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 19.700 7.200 20.950 7.850 ;
        RECT 23.450 7.200 24.050 9.050 ;
        RECT 19.700 7.200 24.050 7.800 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 16.800 8.450 22.700 9.050 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.600 7.800 8.200 9.050 ;
        RECT 2.300 8.450 8.200 9.050 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 25.000 16.250 ;
    END
  END vdd!
  PIN f
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.000 7.200 5.600 7.800 ;
    END
  END f
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.050 10.950 24.500 11.550 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 0.400 4.700 9.550 5.300 ;
        RECT 8.950 4.700 9.550 6.550 ;
        RECT 15.300 5.900 15.900 6.550 ;
        RECT 8.950 5.950 15.900 6.550 ;
        RECT 18.650 5.950 22.700 6.550 ;
        RECT 10.150 4.700 24.400 5.300 ;
  END 
END oai222_4

MACRO oai222_3
  CLASS  CORE ;
  FOREIGN oai222_3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 22.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 10.950 7.200 11.550 9.050 ;
        RECT 10.950 8.450 15.400 9.050 ;
        RECT 14.800 7.700 15.400 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 22.500 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 12.300 7.200 14.300 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 17.200 7.200 18.350 7.800 ;
        RECT 17.650 8.450 21.250 9.050 ;
        RECT 17.650 7.200 18.350 9.050 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 19.650 7.150 20.250 7.800 ;
        RECT 18.850 7.200 20.850 7.800 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.950 7.200 6.550 9.000 ;
        RECT 1.100 8.400 6.550 9.000 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 13.450 13.500 14.150 16.250 ;
        RECT 0.000 13.750 22.500 16.250 ;
    END
  END vdd!
  PIN f
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.000 7.200 4.000 7.800 ;
    END
  END f
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.450 9.700 21.900 10.300 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 0.350 5.950 13.600 6.550 ;
        RECT 16.300 5.950 20.350 6.550 ;
        RECT 11.250 4.700 22.050 5.300 ;
  END 
END oai222_3

MACRO oai222_2
  CLASS  CORE ;
  FOREIGN oai222_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 17.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.550 7.200 8.550 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 17.500 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.050 7.200 11.050 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 11.550 7.200 13.550 7.800 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 14.200 7.200 16.200 7.800 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.700 7.700 5.300 9.050 ;
        RECT 0.950 8.450 5.300 9.050 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 17.500 16.250 ;
    END
  END vdd!
  PIN f
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.100 7.200 4.100 7.800 ;
    END
  END f
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.600 9.700 16.800 10.300 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 2.600 4.700 10.050 5.300 ;
        RECT 7.700 5.900 15.100 6.500 ;
        RECT 12.800 4.700 16.800 5.300 ;
  END 
END oai222_2

MACRO oai222_1
  CLASS  CORE ;
  FOREIGN oai222_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.400 7.200 8.400 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 12.500 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.950 7.200 5.550 8.000 ;
        RECT 3.900 7.200 5.900 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.900 7.200 10.900 7.800 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 10.950 8.450 11.550 10.300 ;
        RECT 10.950 8.450 12.250 9.050 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.300 5.950 2.300 6.550 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 12.500 16.250 ;
    END
  END vdd!
  PIN f
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.500 8.450 3.500 9.050 ;
    END
  END f
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.450 9.700 9.150 10.300 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 2.800 5.950 7.150 6.550 ;
        RECT 2.800 5.950 3.400 7.800 ;
        RECT 2.000 7.200 3.400 7.800 ;
        RECT 8.100 5.950 10.500 6.550 ;
        RECT 4.700 4.700 12.200 5.300 ;
  END 
END oai222_1

MACRO oai221_5
  CLASS  CORE ;
  FOREIGN oai221_5 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 28.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 13.900 8.450 15.900 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 28.750 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 20.850 7.200 22.850 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.200 8.400 5.200 9.050 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 8.450 2.250 9.050 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 24.750 7.200 26.750 7.800 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 5.600 13.550 6.300 16.250 ;
        RECT 0.000 13.750 28.750 16.250 ;
        RECT 25.750 13.500 26.450 16.250 ;
        RECT 21.450 13.550 22.150 16.250 ;
        RECT 16.250 13.550 16.950 16.250 ;
        RECT 10.800 13.550 11.500 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.050 10.950 28.100 11.550 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 3.150 3.450 10.550 4.050 ;
        RECT 11.850 3.450 26.250 4.050 ;
  END 
END oai221_5

MACRO oai221_4
  CLASS  CORE ;
  FOREIGN oai221_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 23.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 14.200 8.350 14.800 9.050 ;
        RECT 14.200 8.450 16.200 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 23.750 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 10.850 8.450 12.850 9.050 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.200 8.450 5.200 9.050 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 8.450 2.250 9.050 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 21.000 8.450 23.000 9.050 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 5.600 13.550 6.300 16.250 ;
        RECT 0.000 13.750 23.750 16.250 ;
        RECT 16.000 13.550 16.700 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.050 10.950 22.650 11.550 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 3.150 3.450 7.250 4.050 ;
        RECT 11.850 3.450 22.650 4.050 ;
  END 
END oai221_4

MACRO oai221_3
  CLASS  CORE ;
  FOREIGN oai221_3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 20.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 17.100 8.450 19.100 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 20.000 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.600 8.450 11.850 9.050 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.200 8.450 5.200 9.050 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.450 7.200 2.450 7.800 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 11.450 7.200 12.200 7.850 ;
        RECT 11.450 7.200 13.450 7.800 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 5.600 13.550 6.300 16.250 ;
        RECT 0.000 13.750 20.000 16.250 ;
        RECT 15.100 13.550 15.800 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.050 10.950 18.400 11.550 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 9.550 4.700 16.950 5.300 ;
        RECT 3.150 3.450 18.650 4.050 ;
  END 
END oai221_3

MACRO oai221_2
  CLASS  CORE ;
  FOREIGN oai221_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.200 7.200 11.200 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 4.800 0.000 5.500 2.700 ;
        RECT 0.000 0.000 15.000 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.700 7.200 8.700 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.500 7.200 3.500 7.800 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.200 7.200 6.200 7.800 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 12.200 7.200 14.200 7.800 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 15.000 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.050 10.950 14.550 11.550 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 3.150 3.450 10.550 4.050 ;
  END 
END oai221_2

MACRO oai221_1
  CLASS  CORE ;
  FOREIGN oai221_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.400 8.400 5.300 9.100 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 11.250 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.900 8.400 7.800 9.100 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.100 5.950 3.100 6.550 ;
        RECT 2.450 5.950 3.100 6.600 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.350 8.450 2.350 9.050 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.400 8.400 10.300 9.100 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 11.250 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.750 4.700 10.750 5.300 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 2.050 4.700 7.350 5.300 ;
  END 
END oai221_1

MACRO oai21_6
  CLASS  CORE ;
  FOREIGN oai21_6 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 17.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.650 7.200 15.400 7.850 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 9.150 0.000 9.850 2.700 ;
        RECT 0.000 0.000 17.500 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.200 5.950 16.050 6.550 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.850 7.200 4.200 7.800 ;
    END
  END c
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 4.050 13.550 4.750 16.250 ;
        RECT 0.000 13.750 17.500 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.400 9.700 16.800 10.300 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 0.700 4.700 11.500 5.300 ;
  END 
END oai21_6

MACRO oai21_5
  CLASS  CORE ;
  FOREIGN oai21_5 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.200 7.200 13.850 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 15.000 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.050 5.950 12.900 6.550 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.850 7.200 2.900 7.800 ;
    END
  END c
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 3.850 13.550 4.450 16.250 ;
        RECT 0.000 13.750 15.000 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.150 9.700 11.950 10.300 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 0.450 4.700 11.250 5.300 ;
  END 
END oai21_5

MACRO oai21_4
  CLASS  CORE ;
  FOREIGN oai21_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.350 7.100 4.950 7.800 ;
        RECT 4.350 7.200 10.400 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 9.850 0.000 10.450 2.550 ;
        RECT 0.000 0.000 12.500 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.950 5.950 12.150 6.550 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 7.200 2.250 7.800 ;
    END
  END c
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 3.650 13.550 4.250 16.250 ;
        RECT 0.000 13.750 12.500 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.950 9.700 12.050 10.300 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 0.350 4.700 12.150 5.300 ;
  END 
END oai21_4

MACRO oai21_3
  CLASS  CORE ;
  FOREIGN oai21_3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.850 5.950 9.750 6.550 ;
        RECT 9.100 5.950 9.750 6.600 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 11.250 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.050 7.200 10.900 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.150 5.950 4.150 6.550 ;
    END
  END c
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 11.250 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.300 9.700 7.950 10.300 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 1.800 3.450 9.200 4.050 ;
  END 
END oai21_3

MACRO oai21_2
  CLASS  CORE ;
  FOREIGN oai21_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.100 5.950 7.000 6.550 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 8.750 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.650 7.200 6.650 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 5.950 2.250 6.550 ;
    END
  END c
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 2.150 13.550 2.750 16.250 ;
        RECT 0.000 13.750 8.750 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.350 9.700 5.400 10.300 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 2.150 4.700 6.150 5.300 ;
  END 
END oai21_2

MACRO oai21_1
  CLASS  CORE ;
  FOREIGN oai21_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.650 8.450 4.650 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 4.250 0.000 4.850 2.600 ;
        RECT 0.000 0.000 7.500 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.450 5.950 6.450 6.550 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.100 5.950 3.100 6.550 ;
    END
  END c
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 7.500 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.850 9.700 5.800 10.300 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 2.550 4.700 6.550 5.300 ;
  END 
END oai21_1

MACRO oai211_5
  CLASS  CORE ;
  FOREIGN oai211_5 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 23.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 21.200 5.950 23.200 6.550 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 23.750 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 12.150 5.950 19.950 6.550 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.050 8.450 4.050 9.050 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.350 8.450 10.400 9.050 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 23.750 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.400 5.950 6.200 6.550 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 2.950 3.450 20.300 4.050 ;
        RECT 2.150 9.700 23.350 10.300 ;
  END 
END oai211_5

MACRO oai211_4
  CLASS  CORE ;
  FOREIGN oai211_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 18.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.300 4.700 9.300 5.300 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 18.750 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.950 7.200 17.900 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.450 8.450 2.450 9.100 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.050 7.200 7.700 7.800 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 18.750 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.950 8.450 11.650 9.050 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 12.550 8.450 16.600 9.050 ;
        RECT 0.300 3.450 16.650 4.050 ;
  END 
END oai211_4

MACRO oai211_3
  CLASS  CORE ;
  FOREIGN oai211_3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 16.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.000 5.950 6.000 6.550 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 16.250 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.500 5.950 9.600 6.550 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 13.400 7.200 15.400 7.800 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 10.400 7.200 12.400 7.800 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 3.800 13.500 4.500 16.250 ;
        RECT 0.000 13.750 16.250 16.250 ;
        RECT 13.400 13.500 14.100 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.000 8.450 15.800 9.050 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 2.150 8.400 6.250 9.000 ;
        RECT 3.100 3.450 15.900 4.050 ;
  END 
END oai211_3

MACRO oai211_2
  CLASS  CORE ;
  FOREIGN oai211_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.350 7.200 9.350 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 12.500 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 10.400 7.200 12.250 7.850 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 7.200 2.250 7.800 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.250 7.200 6.600 7.800 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 12.500 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.300 8.450 6.950 9.050 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 0.300 3.450 10.350 4.050 ;
        RECT 8.050 8.450 12.050 9.050 ;
  END 
END oai211_2

MACRO oai211_1
  CLASS  CORE ;
  FOREIGN oai211_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.850 7.200 3.200 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 10.000 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.350 8.450 5.450 9.050 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.750 7.200 9.750 7.800 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.150 7.200 7.250 7.800 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 10.000 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.000 9.700 9.700 10.300 ;
    END
  END x
END oai211_1

MACRO oa44_6
  CLASS  CORE ;
  FOREIGN oa44_6 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 35.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 27.000 8.450 29.000 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 35.000 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 22.100 8.450 24.100 9.050 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 29.600 7.200 31.600 7.800 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 32.700 7.200 34.700 7.800 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.900 8.450 7.900 9.050 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 35.000 16.250 ;
    END
  END vdd!
  PIN f
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 10.750 8.450 12.750 9.050 ;
    END
  END f
  PIN g
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.400 7.200 5.400 7.800 ;
    END
  END g
  PIN h
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 7.200 2.250 7.800 ;
    END
  END h
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 10.900 7.200 24.000 7.800 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 4.100 3.450 19.600 4.050 ;
        RECT 21.900 3.450 30.800 4.050 ;
  END 
END oa44_6

MACRO oa44_5
  CLASS  CORE ;
  FOREIGN oa44_5 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 33.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 25.850 8.350 27.650 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 9.150 0.000 9.850 2.750 ;
        RECT 0.000 0.000 33.750 2.500 ;
        RECT 23.750 0.000 24.450 2.750 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 22.100 8.350 23.900 9.050 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 28.250 7.200 30.350 7.800 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 31.500 7.200 33.500 7.800 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.850 8.350 7.650 9.050 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 33.750 16.250 ;
    END
  END vdd!
  PIN f
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.700 8.350 10.500 9.050 ;
    END
  END f
  PIN g
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.400 7.200 5.500 7.800 ;
    END
  END g
  PIN h
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 7.200 2.250 7.800 ;
    END
  END h
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 15.850 4.700 17.900 5.300 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 4.100 4.700 12.850 5.300 ;
        RECT 20.450 4.700 29.500 5.300 ;
  END 
END oa44_5

MACRO oa44_4
  CLASS  CORE ;
  FOREIGN oa44_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 25.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 18.350 7.200 21.100 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 4.200 0.000 4.800 2.800 ;
        RECT 0.000 0.000 25.000 2.500 ;
        RECT 20.200 0.000 20.800 2.800 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 17.200 5.950 17.800 7.800 ;
        RECT 15.900 7.200 17.800 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 20.400 5.950 22.400 6.550 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 22.900 5.900 24.750 6.550 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.900 7.200 6.650 7.800 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 25.000 16.250 ;
    END
  END vdd!
  PIN f
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.200 5.950 7.800 7.800 ;
        RECT 7.200 7.200 9.100 7.800 ;
    END
  END f
  PIN g
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.600 5.950 4.600 6.550 ;
    END
  END g
  PIN h
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 5.900 2.100 6.550 ;
    END
  END h
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 10.850 5.950 12.850 6.550 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 2.500 4.700 10.000 5.300 ;
        RECT 9.400 4.700 10.000 5.450 ;
        RECT 15.000 4.700 22.500 5.300 ;
        RECT 15.000 4.700 15.600 5.450 ;
  END 
END oa44_4

MACRO oa44_3
  CLASS  CORE ;
  FOREIGN oa44_3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 25.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 19.600 5.850 21.350 6.550 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 25.000 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 15.850 5.950 17.850 6.550 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 20.400 7.200 22.400 7.800 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 22.900 7.150 24.750 7.800 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.650 5.850 5.400 6.550 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 25.000 16.250 ;
    END
  END vdd!
  PIN f
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.150 5.950 9.150 6.550 ;
    END
  END f
  PIN g
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.600 7.200 4.600 7.800 ;
    END
  END g
  PIN h
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 7.150 2.100 7.800 ;
    END
  END h
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 12.150 4.700 12.850 6.550 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 2.500 4.700 11.150 5.300 ;
        RECT 5.900 4.700 6.500 7.750 ;
        RECT 13.850 4.700 22.500 5.300 ;
        RECT 18.500 4.700 19.100 7.750 ;
  END 
END oa44_3

MACRO oa44_2
  CLASS  CORE ;
  FOREIGN oa44_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 18.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.150 8.100 6.750 9.050 ;
        RECT 4.800 8.350 6.750 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 18.750 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.150 5.950 6.150 6.550 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.650 5.950 3.650 6.550 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.750 8.400 2.750 9.050 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 12.050 8.100 12.650 9.050 ;
        RECT 12.050 8.350 13.850 9.050 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 18.750 16.250 ;
    END
  END vdd!
  PIN f
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 12.650 5.950 14.650 6.550 ;
    END
  END f
  PIN g
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 15.150 5.950 17.150 6.550 ;
    END
  END g
  PIN h
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 15.900 8.400 17.900 9.050 ;
    END
  END h
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.100 5.650 9.700 9.050 ;
        RECT 7.750 8.450 9.700 9.050 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 2.200 4.650 8.600 5.250 ;
        RECT 8.000 4.650 8.600 7.500 ;
        RECT 10.200 4.650 16.600 5.250 ;
        RECT 10.200 4.650 10.800 7.500 ;
  END 
END oa44_2

MACRO oa44_1
  CLASS  CORE ;
  FOREIGN oa44_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 17.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.400 8.450 5.900 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 17.500 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.000 5.950 6.000 6.550 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.500 5.950 3.500 6.550 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.850 8.450 2.850 9.050 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 10.600 8.450 12.600 9.050 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 17.500 16.250 ;
    END
  END vdd!
  PIN f
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 11.500 5.950 13.500 6.550 ;
    END
  END f
  PIN g
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 14.000 5.950 16.000 6.550 ;
    END
  END g
  PIN h
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 15.000 8.450 17.000 9.050 ;
    END
  END h
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.450 7.100 9.050 9.050 ;
        RECT 6.750 8.450 9.050 9.050 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 2.050 4.650 7.500 5.250 ;
        RECT 6.900 4.650 7.500 7.150 ;
        RECT 10.000 4.650 15.900 5.250 ;
        RECT 10.000 4.650 10.600 7.150 ;
  END 
END oa44_1

MACRO oa33_6
  CLASS  CORE ;
  FOREIGN oa33_6 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.400 5.950 2.400 6.550 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 15.000 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.900 5.950 4.900 6.550 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.000 8.450 6.000 9.050 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 11.700 8.400 13.700 9.050 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 10.500 5.850 12.000 6.650 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 15.000 16.250 ;
    END
  END vdd!
  PIN f
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.200 8.400 11.200 9.050 ;
    END
  END f
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.100 5.850 8.850 6.650 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 0.350 4.650 0.950 5.300 ;
        RECT 0.350 4.700 12.850 5.300 ;
        RECT 1.950 7.200 14.550 7.800 ;
        RECT 1.950 7.200 2.550 9.050 ;
  END 
END oa33_6

MACRO oa33_5
  CLASS  CORE ;
  FOREIGN oa33_5 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.750 5.950 7.750 6.550 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 5.700 0.000 6.300 2.950 ;
        RECT 0.000 0.000 13.750 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.250 5.950 5.250 6.550 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.650 8.450 5.650 9.050 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.550 8.300 10.350 9.050 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 10.050 5.950 12.050 6.550 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 13.750 16.250 ;
    END
  END vdd!
  PIN f
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 11.500 8.450 13.500 9.050 ;
    END
  END f
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.400 5.950 2.750 6.550 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 4.000 4.700 11.500 5.300 ;
        RECT 0.850 7.200 13.200 7.800 ;
        RECT 7.400 7.200 8.000 9.200 ;
  END 
END oa33_5

MACRO oa33_4
  CLASS  CORE ;
  FOREIGN oa33_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.400 5.950 6.900 6.750 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 5.700 0.000 6.300 2.950 ;
        RECT 0.000 0.000 13.750 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.250 5.950 4.750 6.750 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.650 8.450 5.650 9.050 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.100 8.450 9.300 9.050 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.450 7.200 11.450 7.800 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 13.750 16.250 ;
    END
  END vdd!
  PIN f
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 11.500 8.450 13.500 9.050 ;
    END
  END f
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.350 5.950 2.750 6.600 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 4.000 3.450 11.500 4.050 ;
        RECT 7.400 5.950 13.200 6.550 ;
        RECT 7.400 5.950 8.000 7.850 ;
        RECT 0.850 7.250 8.000 7.850 ;
  END 
END oa33_4

MACRO oa33_3
  CLASS  CORE ;
  FOREIGN oa33_3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.400 8.450 2.000 9.200 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 2.100 0.000 2.700 3.000 ;
        RECT 0.000 0.000 12.500 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.550 5.950 3.550 6.550 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.600 8.450 4.200 9.200 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 10.250 5.950 12.250 6.550 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.650 8.450 10.650 9.050 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 7.500 13.550 8.100 16.250 ;
        RECT 0.000 13.750 12.500 16.250 ;
    END
  END vdd!
  PIN f
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.750 5.950 9.750 6.550 ;
    END
  END f
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.800 8.450 8.150 9.050 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 7.500 3.300 8.100 4.100 ;
        RECT 0.400 3.500 11.500 4.100 ;
        RECT 4.700 8.450 5.300 10.300 ;
        RECT 0.450 9.700 11.700 10.300 ;
  END 
END oa33_3

MACRO oa33_2
  CLASS  CORE ;
  FOREIGN oa33_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 8.450 2.250 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 1.050 0.000 1.750 2.700 ;
        RECT 0.000 0.000 12.500 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.450 5.950 3.450 6.550 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.750 8.450 4.600 9.100 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 10.250 8.450 12.250 9.050 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.050 5.950 11.050 6.550 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 7.800 13.600 8.500 16.250 ;
        RECT 0.000 13.750 12.500 16.250 ;
    END
  END vdd!
  PIN f
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.600 8.450 9.600 9.050 ;
    END
  END f
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.650 5.950 7.650 6.550 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 2.800 4.700 11.500 5.300 ;
        RECT 5.100 8.450 5.700 10.300 ;
        RECT 0.400 9.700 11.950 10.300 ;
  END 
END oa33_2

MACRO oa33_1
  CLASS  CORE ;
  FOREIGN oa33_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.900 9.700 2.900 10.300 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 11.250 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.700 7.200 2.700 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.400 7.150 5.350 7.850 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.950 7.200 10.950 7.800 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.400 9.700 10.400 10.300 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 4.450 13.550 5.150 16.250 ;
        RECT 0.000 13.750 11.250 16.250 ;
    END
  END vdd!
  PIN f
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.300 7.200 8.300 7.800 ;
    END
  END f
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.850 9.700 7.850 10.300 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 2.750 3.450 10.200 4.050 ;
  END 
END oa33_1

MACRO oa31_6
  CLASS  CORE ;
  FOREIGN oa31_6 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.200 7.100 7.800 9.100 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 11.250 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.450 8.450 6.450 9.050 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.450 5.850 4.150 7.850 ;
        RECT 3.450 5.850 4.650 6.700 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.000 7.200 11.000 7.800 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 11.250 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.950 7.150 1.550 9.150 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 5.150 5.950 9.200 6.550 ;
        RECT 8.450 8.450 10.900 9.050 ;
        RECT 2.200 6.700 2.800 10.300 ;
        RECT 8.450 8.450 9.050 10.300 ;
        RECT 2.200 9.700 9.050 10.300 ;
  END 
END oa31_6

MACRO oa31_5
  CLASS  CORE ;
  FOREIGN oa31_5 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.500 7.200 8.500 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 11.250 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.000 7.200 6.000 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.100 5.950 4.650 6.550 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.000 7.200 11.000 7.800 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 11.250 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.850 8.450 2.900 9.050 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 5.150 5.950 9.200 6.550 ;
        RECT 7.550 8.450 10.950 9.050 ;
  END 
END oa31_5

MACRO oa31_4
  CLASS  CORE ;
  FOREIGN oa31_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.400 7.200 8.400 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 11.250 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.900 7.200 5.900 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.100 5.950 4.650 6.550 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.900 7.200 10.900 7.800 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 11.250 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.850 8.450 2.900 9.050 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 5.150 5.900 9.150 6.500 ;
        RECT 7.500 8.450 10.850 9.050 ;
  END 
END oa31_4

MACRO oa31_3
  CLASS  CORE ;
  FOREIGN oa31_3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.950 7.100 6.550 9.100 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 5.500 0.000 6.200 2.800 ;
        RECT 0.000 0.000 10.000 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.450 7.100 4.050 9.100 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.850 5.950 2.850 6.550 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.550 8.450 9.750 9.050 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 8.350 13.550 9.050 16.250 ;
        RECT 0.000 13.750 10.000 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.400 9.700 7.700 10.300 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 3.800 5.900 7.900 6.500 ;
        RECT 8.950 5.950 9.550 7.800 ;
        RECT 7.200 7.200 9.550 7.800 ;
  END 
END oa31_3

MACRO oa31_2
  CLASS  CORE ;
  FOREIGN oa31_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.950 5.850 6.550 7.900 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 5.400 0.000 6.150 2.650 ;
        RECT 0.000 0.000 8.750 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.400 7.150 5.350 7.850 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.200 4.600 2.800 6.600 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.200 5.850 7.800 7.900 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 8.750 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 7.200 2.250 7.800 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 3.750 4.700 7.750 5.300 ;
  END 
END oa31_2

MACRO oa31_1
  CLASS  CORE ;
  FOREIGN oa31_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.950 5.850 6.550 7.900 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 8.750 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.400 7.150 5.350 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.200 4.600 2.800 6.600 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.200 5.850 7.800 7.900 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 8.750 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 7.200 2.250 7.800 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 3.700 4.700 7.750 5.300 ;
  END 
END oa31_1

MACRO oa22_6
  CLASS  CORE ;
  FOREIGN oa22_6 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.250 7.200 9.150 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.350 0.000 0.950 2.650 ;
        RECT 0.000 0.000 11.250 2.500 ;
        RECT 7.650 0.000 8.350 2.700 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 7.100 1.750 7.900 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.250 5.950 4.250 6.550 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.850 5.950 6.850 6.550 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 6.050 13.500 6.800 16.250 ;
        RECT 0.000 13.750 11.250 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.150 4.700 10.500 5.300 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 2.200 4.700 6.550 5.300 ;
  END 
END oa22_6

MACRO oa22_5
  CLASS  CORE ;
  FOREIGN oa22_5 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.350 7.200 9.150 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 7.150 0.000 7.750 2.700 ;
        RECT 0.000 0.000 11.250 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 7.100 1.750 7.900 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.350 5.950 4.350 6.550 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.850 5.950 6.850 6.550 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 6.100 13.500 6.800 16.250 ;
        RECT 0.000 13.750 11.250 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.350 4.700 10.500 5.300 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 2.050 4.650 6.050 5.250 ;
  END 
END oa22_5

MACRO oa22_4
  CLASS  CORE ;
  FOREIGN oa22_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.900 7.200 6.650 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 7.150 0.000 7.750 2.700 ;
        RECT 0.000 0.000 10.000 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 4.700 2.250 5.300 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.750 4.700 4.750 5.300 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.250 4.700 7.250 5.300 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 10.000 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.450 3.450 9.450 4.050 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 2.050 3.450 6.050 4.050 ;
  END 
END oa22_4

MACRO oa22_3
  CLASS  CORE ;
  FOREIGN oa22_3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.150 5.950 9.150 6.550 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 10.000 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 7.200 2.250 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.750 7.200 4.750 7.800 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.250 7.100 5.850 7.800 ;
        RECT 5.250 7.200 7.250 7.800 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 10.000 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.900 3.450 9.650 4.050 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 2.050 3.450 6.050 4.050 ;
  END 
END oa22_3

MACRO oa22_2
  CLASS  CORE ;
  FOREIGN oa22_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.100 4.700 6.550 5.300 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 10.000 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.950 3.300 1.550 5.300 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.100 5.950 4.150 6.550 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.950 5.950 7.950 6.550 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 5.650 13.550 6.250 16.250 ;
        RECT 0.000 13.750 10.000 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.650 3.450 9.650 4.050 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 2.150 3.450 6.250 4.050 ;
  END 
END oa22_2

MACRO oa22_1
  CLASS  CORE ;
  FOREIGN oa22_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.100 4.700 6.550 5.300 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 10.000 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.950 3.300 1.550 5.300 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.100 5.950 4.100 6.550 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.950 5.950 7.950 6.550 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 10.000 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.650 3.450 9.650 4.050 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 2.150 3.450 6.250 4.050 ;
  END 
END oa22_1

MACRO oa222_5
  CLASS  CORE ;
  FOREIGN oa222_5 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.650 7.100 9.150 7.900 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 5.550 0.000 6.150 2.800 ;
        RECT 0.000 0.000 15.000 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.700 5.850 10.300 7.250 ;
        RECT 9.700 5.850 11.650 6.650 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 13.100 5.850 14.600 6.650 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 11.300 8.350 12.900 9.150 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.650 7.100 7.150 7.900 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 15.000 16.250 ;
    END
  END vdd!
  PIN f
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.300 7.100 4.850 7.900 ;
    END
  END f
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.450 8.450 3.500 9.050 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 3.850 5.800 9.200 6.400 ;
        RECT 7.100 9.700 14.350 10.300 ;
        RECT 6.850 4.700 14.350 5.300 ;
        RECT 11.950 7.200 14.500 7.800 ;
  END 
END oa222_5

MACRO oa222_4
  CLASS  CORE ;
  FOREIGN oa222_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.800 7.100 9.300 7.900 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 5.550 0.000 6.150 2.800 ;
        RECT 0.000 0.000 15.000 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 10.000 5.850 10.750 7.000 ;
        RECT 10.000 5.850 11.650 6.650 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 13.100 5.850 14.600 6.650 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 11.300 8.350 12.900 9.150 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.650 7.100 7.150 7.900 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 15.000 16.250 ;
    END
  END vdd!
  PIN f
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.300 7.100 4.850 7.900 ;
    END
  END f
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.450 8.450 3.500 9.050 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 3.850 5.800 9.200 6.400 ;
        RECT 7.100 9.700 14.350 10.300 ;
        RECT 6.850 4.700 14.350 5.300 ;
        RECT 11.950 7.200 14.500 7.800 ;
  END 
END oa222_4

MACRO oa222_3
  CLASS  CORE ;
  FOREIGN oa222_3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.800 7.100 8.300 7.900 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 13.750 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.800 8.350 10.400 9.150 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 11.450 8.350 12.950 9.150 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 10.850 5.850 11.650 7.750 ;
        RECT 10.200 7.150 11.650 7.750 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.550 7.100 6.300 7.900 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 9.100 13.450 9.700 16.250 ;
        RECT 0.000 13.750 13.750 16.250 ;
    END
  END vdd!
  PIN f
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.100 5.850 3.600 6.650 ;
    END
  END f
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.850 9.700 2.850 10.300 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 3.700 4.700 8.350 5.300 ;
        RECT 5.950 5.900 10.000 6.500 ;
        RECT 6.450 9.700 12.900 10.300 ;
        RECT 11.000 4.750 13.400 5.350 ;
        RECT 12.800 4.750 13.400 6.950 ;
  END 
END oa222_3

MACRO oa222_2
  CLASS  CORE ;
  FOREIGN oa222_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.650 9.700 10.750 10.300 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 5.400 0.000 6.100 2.650 ;
        RECT 0.000 0.000 12.500 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 10.000 7.200 11.950 7.850 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.550 7.200 9.400 7.850 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.950 9.700 6.950 10.300 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.500 5.900 4.250 6.600 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 12.500 16.250 ;
    END
  END vdd!
  PIN f
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.200 9.650 4.100 10.300 ;
    END
  END f
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 5.900 2.000 6.600 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 4.700 7.200 7.050 7.800 ;
        RECT 4.750 5.950 12.200 6.550 ;
  END 
END oa222_2

MACRO oa222_1
  CLASS  CORE ;
  FOREIGN oa222_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.600 9.700 10.600 10.300 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 12.500 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 10.250 7.200 12.250 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.750 7.200 9.750 7.800 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.800 9.700 7.800 10.300 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.400 5.950 4.100 7.800 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 12.500 16.250 ;
    END
  END vdd!
  PIN f
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.950 9.700 2.950 10.300 ;
    END
  END f
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.350 5.950 2.350 6.550 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 4.700 7.200 7.050 7.800 ;
        RECT 4.750 5.950 12.200 6.550 ;
  END 
END oa222_1

MACRO oa221_5
  CLASS  CORE ;
  FOREIGN oa221_5 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.550 8.450 6.550 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 13.750 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.100 7.200 4.300 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.900 7.200 7.950 7.800 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.100 8.450 9.100 9.050 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.350 8.450 2.350 9.050 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 4.000 13.550 4.750 16.250 ;
        RECT 0.000 13.750 13.750 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 11.000 7.200 11.600 10.300 ;
        RECT 11.000 7.200 12.800 7.800 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 3.850 3.450 9.200 4.050 ;
        RECT 9.900 8.500 10.500 10.300 ;
        RECT 0.350 9.700 10.500 10.300 ;
  END 
END oa221_5

MACRO oa221_4
  CLASS  CORE ;
  FOREIGN oa221_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.850 8.450 6.550 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 13.750 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.100 7.200 4.250 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.850 7.200 7.950 7.800 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.100 8.450 9.100 9.050 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 8.450 2.550 9.050 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 13.750 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 11.000 7.200 13.000 7.800 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 3.850 3.450 9.200 4.050 ;
        RECT 9.900 6.900 10.500 10.300 ;
        RECT 0.350 9.700 10.500 10.300 ;
  END 
END oa221_4

MACRO oa221_3
  CLASS  CORE ;
  FOREIGN oa221_3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.850 8.450 6.500 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 13.750 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.100 7.200 4.250 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.850 7.200 8.000 7.800 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.150 8.450 9.150 9.050 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 8.450 2.550 9.050 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 13.750 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 11.100 7.200 13.100 7.800 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 3.850 3.450 9.200 4.050 ;
        RECT 9.800 7.950 10.400 10.300 ;
        RECT 0.350 9.700 10.400 10.300 ;
  END 
END oa221_3

MACRO oa221_2
  CLASS  CORE ;
  FOREIGN oa221_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.850 8.450 6.000 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 11.250 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.100 7.200 4.250 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.650 7.200 7.700 7.800 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.500 8.450 8.500 9.050 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 8.450 2.550 9.050 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 7.900 13.500 8.600 16.250 ;
        RECT 0.000 13.750 11.250 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.500 7.200 10.900 7.800 ;
        RECT 10.300 7.200 10.900 8.000 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 8.500 3.000 9.100 4.050 ;
        RECT 3.850 3.450 9.100 4.050 ;
        RECT 9.150 8.400 9.750 10.300 ;
        RECT 1.050 9.700 9.750 10.300 ;
  END 
END oa221_2

MACRO oa221_1
  CLASS  CORE ;
  FOREIGN oa221_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.300 8.450 5.300 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 10.000 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.350 7.200 3.350 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.850 7.200 7.850 7.800 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.650 8.450 9.750 9.050 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 8.450 2.250 9.050 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 10.000 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.100 3.450 9.550 4.050 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 0.350 9.700 5.250 10.300 ;
        RECT 2.150 4.700 6.150 5.300 ;
  END 
END oa221_1

MACRO oa21_6
  CLASS  CORE ;
  FOREIGN oa21_6 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.450 5.950 4.050 6.550 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 6.850 0.000 7.450 2.800 ;
        RECT 0.000 0.000 10.000 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.800 7.200 5.900 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.950 7.500 1.550 9.050 ;
        RECT 0.250 8.450 1.550 9.050 ;
    END
  END c
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 10.000 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.600 5.950 9.600 6.550 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 0.350 3.450 5.750 4.050 ;
        RECT 2.150 8.500 8.400 9.100 ;
  END 
END oa21_6

MACRO oa21_5
  CLASS  CORE ;
  FOREIGN oa21_5 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.900 5.950 3.950 6.550 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 10.000 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.900 7.200 6.000 7.850 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.950 7.500 1.550 9.050 ;
        RECT 0.250 8.450 1.550 9.050 ;
    END
  END c
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.450 13.450 1.050 16.250 ;
        RECT 0.000 13.750 10.000 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.600 5.950 9.600 6.550 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 0.350 4.700 5.750 5.300 ;
        RECT 2.150 8.500 5.850 9.100 ;
  END 
END oa21_5

MACRO oa21_4
  CLASS  CORE ;
  FOREIGN oa21_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.150 5.650 3.750 6.600 ;
        RECT 2.200 5.850 3.750 6.600 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 8.750 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.300 5.850 6.000 6.600 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.950 7.650 1.550 9.050 ;
        RECT 0.300 8.450 1.550 9.050 ;
    END
  END c
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.450 13.450 1.050 16.250 ;
        RECT 0.000 13.750 8.750 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.500 5.950 8.500 6.550 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 2.050 4.550 4.850 5.150 ;
        RECT 4.250 4.550 4.850 5.250 ;
        RECT 0.350 4.700 2.650 5.300 ;
        RECT 2.150 8.500 5.450 9.100 ;
  END 
END oa21_4

MACRO oa21_3
  CLASS  CORE ;
  FOREIGN oa21_3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.100 5.950 4.100 6.550 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 8.750 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.500 7.200 6.500 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.950 7.450 1.550 9.050 ;
        RECT 0.500 8.450 1.550 9.050 ;
    END
  END c
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 8.750 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.450 5.950 8.450 6.550 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 0.350 4.700 4.850 5.300 ;
        RECT 2.150 8.500 6.350 9.100 ;
  END 
END oa21_3

MACRO oa21_2
  CLASS  CORE ;
  FOREIGN oa21_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.000 5.950 4.050 6.550 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 1.400 0.000 2.100 2.950 ;
        RECT 0.000 0.000 7.500 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.650 5.950 6.550 6.600 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.600 7.200 2.600 7.800 ;
    END
  END c
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.450 13.450 1.050 16.250 ;
        RECT 0.000 13.750 7.500 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.150 7.200 7.150 7.800 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 0.450 3.450 3.750 4.050 ;
        RECT 0.450 3.450 1.050 6.200 ;
        RECT 2.150 8.500 5.350 9.100 ;
  END 
END oa21_2

MACRO oa21_1
  CLASS  CORE ;
  FOREIGN oa21_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.300 4.700 2.300 5.300 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 7.500 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.250 8.450 7.250 9.050 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.150 7.200 3.150 7.800 ;
    END
  END c
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 7.500 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.150 5.950 6.150 6.550 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 1.000 8.450 4.750 9.050 ;
  END 
END oa21_1

MACRO oa211_5
  CLASS  CORE ;
  FOREIGN oa211_5 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.100 7.150 9.950 7.850 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 12.500 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 10.450 7.150 12.200 7.850 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.300 7.200 7.600 7.800 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.800 7.200 4.800 7.800 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 4.550 13.500 5.250 16.250 ;
        RECT 0.000 13.750 12.500 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.300 7.200 2.300 7.800 ;
    END
  END x
END oa211_5

MACRO oa211_4
  CLASS  CORE ;
  FOREIGN oa211_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.100 7.200 10.000 7.850 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 12.500 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 10.500 7.150 12.250 7.850 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.600 7.200 7.600 7.800 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.900 7.200 4.900 7.800 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 12.500 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.400 7.200 2.400 7.800 ;
    END
  END x
END oa211_4

MACRO oa211_3
  CLASS  CORE ;
  FOREIGN oa211_3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.750 7.150 8.500 7.850 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 11.250 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.000 7.200 11.000 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.250 7.200 6.250 7.800 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.600 7.200 3.600 7.800 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 3.800 13.500 4.500 16.250 ;
        RECT 0.000 13.750 11.250 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.300 9.700 2.300 10.300 ;
    END
  END x
END oa211_3

MACRO oa211_2
  CLASS  CORE ;
  FOREIGN oa211_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.850 5.950 7.850 6.550 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 8.750 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.500 8.450 8.500 9.050 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.550 8.450 4.600 9.050 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.450 7.150 4.150 7.800 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 8.750 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.350 4.700 2.400 5.300 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 0.350 5.950 5.350 6.550 ;
        RECT 4.750 5.950 5.350 7.800 ;
        RECT 0.350 5.950 0.950 9.050 ;
        RECT 0.350 8.450 2.050 9.050 ;
        RECT 5.100 7.200 5.700 9.050 ;
        RECT 4.350 4.700 8.350 5.300 ;
  END 
END oa211_2

MACRO oa211_1
  CLASS  CORE ;
  FOREIGN oa211_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.900 8.450 7.900 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 8.750 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.450 5.950 8.450 6.550 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.800 8.450 4.800 9.050 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.050 5.950 4.050 6.550 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 8.750 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.300 8.450 2.300 9.050 ;
    END
  END x
END oa211_1

MACRO nor3i_5
  CLASS  CORE ;
  FOREIGN nor3i_5 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 18.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.700 4.700 6.750 5.300 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 18.750 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 12.300 5.950 14.300 6.550 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 15.750 5.950 17.750 6.550 ;
    END
  END c
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 1.750 13.550 2.350 16.250 ;
        RECT 0.000 13.750 18.750 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.200 3.450 18.400 4.050 ;
    END
  END x
END nor3i_5

MACRO nor3i_4
  CLASS  CORE ;
  FOREIGN nor3i_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 16.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.250 3.450 4.250 4.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 16.250 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.800 4.700 11.800 5.300 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 13.250 5.950 15.250 6.550 ;
    END
  END c
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 16.250 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.700 3.450 15.900 4.050 ;
    END
  END x
END nor3i_4

MACRO nor3i_3
  CLASS  CORE ;
  FOREIGN nor3i_3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.800 4.700 2.800 5.300 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 13.750 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.750 6.700 8.350 7.800 ;
        RECT 7.200 7.200 13.300 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.550 5.950 11.550 6.550 ;
    END
  END c
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 5.500 13.550 6.200 16.250 ;
        RECT 0.000 13.750 13.750 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.600 4.700 11.600 5.300 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 4.100 5.750 4.700 6.550 ;
        RECT 0.450 5.950 4.700 6.550 ;
        RECT 3.850 8.450 13.350 9.050 ;
  END 
END nor3i_3

MACRO nor3i_2
  CLASS  CORE ;
  FOREIGN nor3i_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.900 4.700 3.000 5.300 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 11.250 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.200 7.200 9.200 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.700 5.950 7.950 6.550 ;
    END
  END c
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 2.400 13.550 3.100 16.250 ;
        RECT 0.000 13.750 11.250 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.050 4.700 10.150 5.300 ;
    END
  END x
END nor3i_2

MACRO nor3i_1
  CLASS  CORE ;
  FOREIGN nor3i_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.850 7.200 2.850 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 7.500 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.050 5.950 4.550 6.550 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.250 4.700 5.950 5.450 ;
        RECT 5.250 4.700 7.250 5.300 ;
    END
  END c
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 7.500 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.400 3.350 4.050 4.050 ;
        RECT 3.400 3.450 7.150 4.050 ;
    END
  END x
END nor3i_1

MACRO nor3i_0
  CLASS  CORE ;
  FOREIGN nor3i_0 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.850 7.200 2.850 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 7.500 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.350 5.950 5.350 6.550 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.000 4.700 7.050 5.300 ;
    END
  END c
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 7.500 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.400 3.450 7.150 4.050 ;
    END
  END x
END nor3i_0

MACRO nor3_5
  CLASS  CORE ;
  FOREIGN nor3_5 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 16.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.600 5.950 15.450 6.550 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 16.250 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.600 7.200 15.500 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.850 8.450 2.900 9.050 ;
    END
  END c
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 7.800 13.550 8.500 16.250 ;
        RECT 0.000 13.750 16.250 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.400 3.450 10.300 4.050 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 4.200 8.450 12.100 9.050 ;
  END 
END nor3_5

MACRO nor3_4
  CLASS  CORE ;
  FOREIGN nor3_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.450 5.950 12.050 6.550 ;
        RECT 11.350 5.950 12.050 7.850 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 3.750 0.000 4.350 2.700 ;
        RECT 0.000 0.000 13.750 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.200 7.200 10.200 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.950 8.450 2.950 9.050 ;
    END
  END c
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 8.600 13.550 9.200 16.250 ;
        RECT 0.000 13.750 13.750 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.100 8.450 13.400 9.050 ;
    END
  END x
END nor3_4

MACRO nor3_3
  CLASS  CORE ;
  FOREIGN nor3_3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.000 5.950 10.450 6.550 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 4.050 0.000 4.750 2.700 ;
        RECT 0.000 0.000 12.500 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.550 7.200 3.650 7.800 ;
        RECT 5.250 7.200 9.100 7.800 ;
        RECT 2.450 7.300 5.900 7.900 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.050 8.450 7.800 9.050 ;
    END
  END c
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 12.500 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.150 5.950 4.750 6.800 ;
        RECT 4.700 4.700 11.750 5.300 ;
        RECT 2.300 5.950 5.300 6.550 ;
        RECT 4.700 4.700 5.300 6.550 ;
    END
  END x
END nor3_3

MACRO nor3_2
  CLASS  CORE ;
  FOREIGN nor3_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.100 5.900 7.050 6.550 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 8.750 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.950 7.200 6.500 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.850 8.450 7.800 9.050 ;
        RECT 7.200 8.450 7.800 9.100 ;
    END
  END c
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 8.750 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.950 4.700 4.600 6.550 ;
        RECT 3.950 4.700 6.300 5.300 ;
        RECT 2.100 5.950 4.600 6.550 ;
    END
  END x
END nor3_2

MACRO nor3_1
  CLASS  CORE ;
  FOREIGN nor3_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.750 5.950 5.750 6.550 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 6.250 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.200 5.950 3.200 6.550 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.850 8.450 2.850 9.050 ;
    END
  END c
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 6.250 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.850 3.450 5.900 4.050 ;
    END
  END x
END nor3_1

MACRO nor3_0
  CLASS  CORE ;
  FOREIGN nor3_0 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.750 8.450 5.750 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 6.250 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.300 5.950 5.300 6.550 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.850 8.450 2.850 9.050 ;
    END
  END c
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 6.250 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.850 3.450 5.900 4.050 ;
    END
  END x
END nor3_0

MACRO nor2i_8
  CLASS  CORE ;
  FOREIGN nor2i_8 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 16.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.850 7.200 15.850 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 16.250 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 13.900 3.450 15.900 4.050 ;
    END
  END b
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 9.450 13.550 10.150 16.250 ;
        RECT 0.000 13.750 16.250 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.850 9.700 12.750 10.300 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 9.100 3.450 13.100 4.050 ;
  END 
END nor2i_8

MACRO nor2i_6
  CLASS  CORE ;
  FOREIGN nor2i_6 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.700 5.950 2.700 6.550 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 13.750 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.250 4.700 10.250 5.300 ;
    END
  END b
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 9.800 13.550 10.400 16.250 ;
        RECT 0.000 13.750 13.750 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.400 3.450 11.550 4.050 ;
        RECT 7.000 5.950 12.100 6.550 ;
        RECT 10.950 3.450 11.550 6.550 ;
    END
  END x
END nor2i_6

MACRO nor2i_5
  CLASS  CORE ;
  FOREIGN nor2i_5 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.550 7.200 2.550 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 13.750 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.900 7.200 9.900 7.800 ;
    END
  END b
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 9.600 13.550 10.300 16.250 ;
        RECT 0.000 13.750 13.750 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.850 9.700 13.050 10.300 ;
    END
  END x
END nor2i_5

MACRO nor2i_4
  CLASS  CORE ;
  FOREIGN nor2i_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.500 5.950 2.500 6.550 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 3.150 0.000 3.850 2.700 ;
        RECT 0.000 0.000 11.250 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.750 5.950 6.750 6.550 ;
    END
  END b
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 2.100 13.550 2.800 16.250 ;
        RECT 0.000 13.750 11.250 16.250 ;
        RECT 7.550 13.550 8.250 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.700 8.450 10.800 9.050 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 0.450 8.450 4.100 9.050 ;
  END 
END nor2i_4

MACRO nor2i_3
  CLASS  CORE ;
  FOREIGN nor2i_3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.550 5.950 2.550 6.550 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 3.200 0.000 3.800 2.700 ;
        RECT 0.000 0.000 8.750 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.250 5.950 7.250 6.550 ;
    END
  END b
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 2.100 13.550 2.800 16.250 ;
        RECT 0.000 13.750 8.750 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.600 8.450 5.600 9.050 ;
    END
  END x
END nor2i_3

MACRO nor2i_2
  CLASS  CORE ;
  FOREIGN nor2i_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.500 7.200 2.500 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 3.200 0.000 3.800 2.700 ;
        RECT 0.000 0.000 8.750 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.750 7.200 6.750 7.800 ;
    END
  END b
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 2.150 13.550 2.750 16.250 ;
        RECT 0.000 13.750 8.750 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.600 9.700 5.600 10.300 ;
    END
  END x
END nor2i_2

MACRO nor2i_1
  CLASS  CORE ;
  FOREIGN nor2i_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 8.450 2.250 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 1.800 0.000 2.400 2.700 ;
        RECT 0.000 0.000 6.250 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.400 8.450 5.500 9.050 ;
    END
  END b
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 2.150 13.550 2.750 16.250 ;
        RECT 0.000 13.750 6.250 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.450 5.950 5.800 6.550 ;
        RECT 5.200 5.950 5.800 7.850 ;
    END
  END x
END nor2i_1

MACRO nor2i_0
  CLASS  CORE ;
  FOREIGN nor2i_0 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 8.450 2.250 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 6.250 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.900 8.450 5.900 9.050 ;
    END
  END b
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 6.250 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.450 5.950 5.800 6.550 ;
        RECT 5.200 5.950 5.800 7.850 ;
    END
  END x
END nor2i_0

MACRO nor2_8
  CLASS  CORE ;
  FOREIGN nor2_8 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.400 7.200 3.400 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 15.000 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.400 4.700 2.400 5.300 ;
    END
  END b
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 15.000 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.150 4.700 14.650 5.300 ;
    END
  END x
END nor2_8

MACRO nor2_6
  CLASS  CORE ;
  FOREIGN nor2_6 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.400 7.200 3.400 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 12.500 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.400 4.700 2.600 5.300 ;
    END
  END b
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 12.500 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.150 4.700 12.150 5.300 ;
    END
  END x
END nor2_6

MACRO nor2_5
  CLASS  CORE ;
  FOREIGN nor2_5 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.900 7.200 2.900 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 11.250 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.400 4.700 2.400 5.300 ;
    END
  END b
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 11.250 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.800 4.700 10.900 5.300 ;
    END
  END x
END nor2_5

MACRO nor2_4
  CLASS  CORE ;
  FOREIGN nor2_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.600 5.950 9.600 6.550 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 10.000 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.350 4.700 3.350 5.300 ;
    END
  END b
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 10.000 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.500 9.700 8.500 10.300 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 1.850 12.350 9.250 12.950 ;
  END 
END nor2_4

MACRO nor2_3
  CLASS  CORE ;
  FOREIGN nor2_3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.450 7.200 8.450 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 8.750 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.650 7.200 2.650 7.800 ;
    END
  END b
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 8.750 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.150 9.700 8.200 10.300 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 2.450 12.500 6.500 13.100 ;
  END 
END nor2_3

MACRO nor2_2
  CLASS  CORE ;
  FOREIGN nor2_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.100 5.950 7.100 6.550 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 7.500 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.650 5.950 2.650 6.550 ;
    END
  END b
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 7.500 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.350 7.200 5.350 7.800 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 2.450 9.700 6.500 10.300 ;
  END 
END nor2_2

MACRO nor2_1
  CLASS  CORE ;
  FOREIGN nor2_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.750 4.700 4.750 5.300 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 5.000 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 8.450 2.300 9.050 ;
    END
  END b
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 5.000 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.200 7.200 4.550 7.800 ;
    END
  END x
END nor2_1

MACRO nor2_0
  CLASS  CORE ;
  FOREIGN nor2_0 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.250 4.700 4.250 5.300 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 5.000 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 8.450 2.250 9.050 ;
    END
  END b
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 5.000 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.150 7.200 4.550 7.800 ;
    END
  END x
END nor2_0

MACRO nand4i_5
  CLASS  CORE ;
  FOREIGN nand4i_5 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 25.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 22.050 7.200 24.100 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 23.350 0.000 23.950 2.700 ;
        RECT 0.000 0.000 25.000 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 15.900 7.200 19.050 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.900 8.450 8.550 9.050 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 8.450 2.250 9.050 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 2.400 13.550 3.100 16.250 ;
        RECT 0.000 13.750 25.000 16.250 ;
        RECT 12.650 13.550 13.350 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.750 10.950 18.450 11.550 ;
    END
  END x
END nand4i_5

MACRO nand4i_4
  CLASS  CORE ;
  FOREIGN nand4i_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 21.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 18.850 8.450 20.850 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 3.600 0.000 4.200 2.650 ;
        RECT 0.000 0.000 21.250 2.500 ;
        RECT 13.200 0.000 13.800 2.650 ;
        RECT 11.950 0.000 12.550 2.650 ;
        RECT 10.500 0.000 11.100 2.650 ;
        RECT 9.150 0.000 9.750 2.650 ;
        RECT 7.900 0.000 8.500 2.650 ;
        RECT 6.400 0.000 7.000 2.650 ;
        RECT 4.900 0.000 5.500 2.650 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 11.700 8.450 13.700 9.050 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.350 8.450 6.350 9.050 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 8.450 2.250 9.050 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 21.250 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.450 10.950 14.700 11.550 ;
    END
  END x
END nand4i_4

MACRO nand4i_3
  CLASS  CORE ;
  FOREIGN nand4i_3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 17.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.750 8.450 2.750 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 17.500 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.850 7.200 7.850 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 11.250 7.200 13.250 7.800 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 14.600 8.450 16.600 9.050 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 10.850 13.500 11.450 16.250 ;
        RECT 0.000 13.750 17.500 16.250 ;
        RECT 14.300 13.550 14.900 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.750 9.700 16.600 10.300 ;
    END
  END x
END nand4i_3

MACRO nand4i_2
  CLASS  CORE ;
  FOREIGN nand4i_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.750 8.450 2.750 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 15.000 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.900 7.200 6.950 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.350 7.200 11.350 7.800 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 11.900 8.450 14.150 9.050 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 15.000 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.550 9.700 12.950 10.300 ;
    END
  END x
END nand4i_2

MACRO nand4i_1
  CLASS  CORE ;
  FOREIGN nand4i_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 7.200 2.250 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 2.050 0.000 2.650 2.700 ;
        RECT 0.000 0.000 10.000 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.750 7.200 9.750 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.950 7.200 6.600 9.100 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.000 7.900 4.600 9.050 ;
        RECT 2.650 8.450 4.600 9.050 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 2.150 13.550 2.750 16.250 ;
        RECT 0.000 13.750 10.000 16.250 ;
        RECT 8.950 13.650 9.550 16.250 ;
        RECT 5.550 13.550 6.150 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.050 8.450 9.650 10.300 ;
        RECT 3.850 9.700 9.650 10.300 ;
    END
  END x
END nand4i_1

MACRO nand4_5
  CLASS  CORE ;
  FOREIGN nand4_5 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 22.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 17.200 7.200 19.850 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 22.500 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 19.350 9.700 21.350 10.300 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 19.850 12.200 21.900 12.800 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.350 4.600 2.600 5.400 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 18.150 9.600 18.750 16.250 ;
        RECT 0.000 13.750 22.500 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.000 7.200 4.100 7.800 ;
    END
  END x
END nand4_5

MACRO nand4_4
  CLASS  CORE ;
  FOREIGN nand4_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 18.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.450 7.200 2.450 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 17.800 0.000 18.400 3.450 ;
        RECT 0.000 0.000 18.750 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.300 7.200 11.300 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 13.000 8.450 15.000 9.050 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 16.250 7.200 18.300 7.800 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 10.850 13.550 11.550 16.250 ;
        RECT 0.000 13.750 18.750 16.250 ;
        RECT 14.250 13.550 14.950 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.350 10.950 16.600 11.550 ;
    END
  END x
END nand4_4

MACRO nand4_3
  CLASS  CORE ;
  FOREIGN nand4_3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 16.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.450 7.200 2.450 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 15.300 0.000 15.900 3.450 ;
        RECT 0.000 0.000 16.250 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.800 7.200 7.800 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.500 8.450 11.500 9.050 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 13.500 7.200 15.300 7.800 ;
        RECT 14.700 7.200 15.300 8.300 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 7.300 13.550 8.000 16.250 ;
        RECT 0.000 13.750 16.250 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.250 9.700 13.050 10.300 ;
    END
  END x
END nand4_3

MACRO nand4_2
  CLASS  CORE ;
  FOREIGN nand4_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.650 7.200 2.650 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 12.800 0.000 13.400 3.500 ;
        RECT 0.000 0.000 13.750 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.100 7.200 7.100 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.450 8.000 9.050 9.050 ;
        RECT 7.900 8.450 9.750 9.050 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 11.200 8.450 13.200 9.050 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 13.750 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.650 9.700 11.450 10.300 ;
    END
  END x
END nand4_2

MACRO nand4_1
  CLASS  CORE ;
  FOREIGN nand4_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.100 7.200 8.100 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 2.100 0.000 2.700 2.700 ;
        RECT 0.000 0.000 8.750 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.550 7.200 5.550 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.650 5.950 3.000 6.550 ;
        RECT 2.300 5.950 3.000 8.900 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.950 7.150 1.550 9.050 ;
        RECT 0.950 8.450 1.800 9.050 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 7.300 13.600 7.900 16.250 ;
        RECT 0.000 13.750 8.750 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.500 8.450 8.100 10.300 ;
        RECT 2.150 9.700 8.100 10.300 ;
    END
  END x
END nand4_1

MACRO nand3i_5
  CLASS  CORE ;
  FOREIGN nand3i_5 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 16.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.900 7.200 4.700 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 4.400 0.000 5.150 2.700 ;
        RECT 0.000 0.000 16.250 2.500 ;
        RECT 11.600 0.000 12.300 2.700 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.950 5.950 12.300 6.550 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.050 7.200 14.750 7.800 ;
    END
  END c
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 16.250 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.500 9.700 14.100 10.300 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 8.150 4.700 15.900 5.300 ;
  END 
END nand3i_5

MACRO nand3i_4
  CLASS  CORE ;
  FOREIGN nand3i_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.350 7.200 2.550 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 9.800 0.000 10.500 2.700 ;
        RECT 0.000 0.000 15.000 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 11.550 5.950 13.550 6.550 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.600 7.200 13.450 7.800 ;
    END
  END c
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 15.000 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.750 8.450 14.650 9.050 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 0.350 5.950 9.550 6.550 ;
        RECT 3.050 5.950 3.650 6.950 ;
  END 
END nand3i_4

MACRO nand3i_3
  CLASS  CORE ;
  FOREIGN nand3i_3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.550 7.200 2.800 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 11.250 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.350 5.950 8.850 6.550 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.950 7.200 10.250 7.800 ;
        RECT 9.650 7.200 10.250 7.900 ;
    END
  END c
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 11.250 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.200 8.450 8.500 9.050 ;
    END
  END x
END nand3i_3

MACRO nand3i_2
  CLASS  CORE ;
  FOREIGN nand3i_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.550 7.200 3.250 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 8.750 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.350 8.450 5.750 9.050 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.400 8.450 8.450 9.050 ;
    END
  END c
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 8.750 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.300 9.700 8.500 10.300 ;
    END
  END x
END nand3i_2

MACRO nand3i_1
  CLASS  CORE ;
  FOREIGN nand3i_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.850 8.450 2.850 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 7.500 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.200 7.200 5.200 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.600 8.450 6.650 9.050 ;
    END
  END c
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 7.500 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.450 9.700 7.150 10.300 ;
    END
  END x
END nand3i_1

MACRO nand3i_0
  CLASS  CORE ;
  FOREIGN nand3i_0 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.850 8.450 2.850 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 7.500 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.200 7.200 5.200 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.600 5.950 6.650 6.550 ;
    END
  END c
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 7.500 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.400 9.700 7.150 10.300 ;
    END
  END x
END nand3i_0

MACRO nand3_5
  CLASS  CORE ;
  FOREIGN nand3_5 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.450 7.200 5.450 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.300 0.000 1.000 3.550 ;
        RECT 0.000 0.000 13.750 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.950 7.200 11.950 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.350 7.200 2.350 7.800 ;
    END
  END c
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 13.750 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.600 9.700 11.400 10.300 ;
    END
  END x
END nand3_5

MACRO nand3_4
  CLASS  CORE ;
  FOREIGN nand3_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.350 7.200 2.350 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 12.500 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.250 5.950 6.250 6.550 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.100 7.200 11.100 7.800 ;
    END
  END c
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 4.100 13.500 4.800 16.250 ;
        RECT 0.000 13.750 12.500 16.250 ;
        RECT 7.500 13.500 8.200 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.450 9.700 9.850 10.300 ;
    END
  END x
END nand3_4

MACRO nand3_3
  CLASS  CORE ;
  FOREIGN nand3_3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.350 7.200 2.350 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 10.000 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.950 7.200 6.600 9.100 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.150 7.200 9.150 7.800 ;
    END
  END c
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 10.000 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.450 9.700 7.850 10.300 ;
    END
  END x
END nand3_3

MACRO nand3_2
  CLASS  CORE ;
  FOREIGN nand3_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.000 7.200 7.000 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 10.000 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.300 7.200 3.300 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.650 7.200 9.650 7.800 ;
    END
  END c
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 10.000 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.450 9.700 7.850 10.300 ;
    END
  END x
END nand3_2

MACRO nand3_1
  CLASS  CORE ;
  FOREIGN nand3_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.450 8.450 2.450 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 6.250 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.400 7.200 4.050 9.100 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.700 8.450 5.300 10.450 ;
    END
  END c
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 6.250 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.450 9.700 4.100 10.300 ;
        RECT 3.500 9.700 4.100 10.900 ;
    END
  END x
END nand3_1

MACRO nand2i_8
  CLASS  CORE ;
  FOREIGN nand2i_8 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 20.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 17.000 8.450 19.000 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 4.000 0.000 4.700 2.700 ;
        RECT 0.000 0.000 20.000 2.500 ;
        RECT 9.200 0.000 9.900 2.700 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.700 5.950 11.200 6.550 ;
    END
  END b
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 20.000 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.550 7.200 15.100 7.800 ;
    END
  END x
END nand2i_8

MACRO nand2i_6
  CLASS  CORE ;
  FOREIGN nand2i_6 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 16.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 12.750 7.200 14.750 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 16.250 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.850 7.200 2.900 7.800 ;
    END
  END b
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 16.250 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.650 5.950 7.800 6.550 ;
        RECT 2.550 8.450 10.050 9.050 ;
        RECT 7.200 5.950 7.800 9.050 ;
    END
  END x
END nand2i_6

MACRO nand2i_5
  CLASS  CORE ;
  FOREIGN nand2i_5 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.850 8.450 3.000 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 13.750 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.300 7.200 11.350 7.800 ;
    END
  END b
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 13.750 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.550 9.700 13.100 10.300 ;
    END
  END x
END nand2i_5

MACRO nand2i_4
  CLASS  CORE ;
  FOREIGN nand2i_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.850 5.950 10.850 6.550 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 3.800 0.000 4.500 2.750 ;
        RECT 0.000 0.000 12.500 2.500 ;
        RECT 9.100 0.000 9.800 2.750 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.100 7.200 4.600 7.800 ;
    END
  END b
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 12.500 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.350 8.450 6.450 9.050 ;
    END
  END x
END nand2i_4

MACRO nand2i_3
  CLASS  CORE ;
  FOREIGN nand2i_3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.350 7.200 3.350 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 3.150 0.000 3.850 2.700 ;
        RECT 0.000 0.000 8.750 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.400 4.700 8.400 5.300 ;
    END
  END b
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 8.750 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.050 9.700 8.500 10.300 ;
    END
  END x
END nand2i_3

MACRO nand2i_2
  CLASS  CORE ;
  FOREIGN nand2i_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 7.200 2.450 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 6.250 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.150 7.200 5.150 7.800 ;
    END
  END b
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 6.250 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.500 8.450 5.850 9.050 ;
    END
  END x
END nand2i_2

MACRO nand2i_1
  CLASS  CORE ;
  FOREIGN nand2i_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.850 9.700 2.850 10.300 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 6.250 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.900 7.200 3.900 7.800 ;
    END
  END b
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 6.250 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.500 8.450 5.850 9.050 ;
    END
  END x
END nand2i_1

MACRO nand2i_0
  CLASS  CORE ;
  FOREIGN nand2i_0 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.850 9.700 2.850 10.300 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 6.250 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.900 7.200 3.900 7.800 ;
    END
  END b
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 6.250 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.500 8.450 5.850 9.050 ;
    END
  END x
END nand2i_0

MACRO nand3_0
  CLASS  CORE ;
  FOREIGN nand3_0 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.450 8.450 2.450 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 6.250 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.150 7.200 4.150 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.950 8.450 5.950 9.050 ;
    END
  END c
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 6.250 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.350 9.700 4.100 10.300 ;
    END
  END x
END nand3_0

MACRO nand2_8
  CLASS  CORE ;
  FOREIGN nand2_8 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.800 7.200 7.900 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 6.750 0.000 7.350 2.700 ;
        RECT 0.000 0.000 12.500 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.850 7.200 2.850 7.800 ;
    END
  END b
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 12.500 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.100 9.700 10.400 10.300 ;
    END
  END x
END nand2_8

MACRO nand2_6
  CLASS  CORE ;
  FOREIGN nand2_6 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.850 7.200 7.900 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 10.000 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.850 7.200 2.850 7.800 ;
    END
  END b
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 10.000 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.100 9.700 9.650 10.300 ;
    END
  END x
END nand2_6

MACRO nand2_5
  CLASS  CORE ;
  FOREIGN nand2_5 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.850 7.200 7.900 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 8.750 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.950 7.200 1.550 9.200 ;
    END
  END b
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 8.750 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.150 9.700 6.650 10.300 ;
    END
  END x
END nand2_5

MACRO nand2_4
  CLASS  CORE ;
  FOREIGN nand2_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.500 7.200 6.500 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 2.700 0.000 3.300 2.700 ;
        RECT 0.000 0.000 8.750 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.000 7.200 4.000 7.800 ;
    END
  END b
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 8.750 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.300 9.700 6.650 10.300 ;
    END
  END x
END nand2_4

MACRO nand2_3
  CLASS  CORE ;
  FOREIGN nand2_3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.950 7.200 5.950 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 7.500 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.450 7.200 3.450 7.800 ;
    END
  END b
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 4.550 13.550 5.150 16.250 ;
        RECT 0.000 13.750 7.500 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.750 9.700 6.950 10.300 ;
    END
  END x
END nand2_3

MACRO nand2_2
  CLASS  CORE ;
  FOREIGN nand2_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.750 7.200 4.750 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 5.000 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 7.200 2.250 7.800 ;
    END
  END b
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 5.000 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.200 8.450 2.800 10.300 ;
        RECT 2.200 8.450 4.650 9.050 ;
    END
  END x
END nand2_2

MACRO nand2_1
  CLASS  CORE ;
  FOREIGN nand2_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.750 5.950 4.750 6.550 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 5.000 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 5.950 2.250 6.550 ;
    END
  END b
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 5.000 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.100 8.450 4.650 9.050 ;
    END
  END x
END nand2_1

MACRO nand2_0
  CLASS  CORE ;
  FOREIGN nand2_0 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.750 7.200 4.750 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 5.000 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 7.200 2.250 7.800 ;
    END
  END b
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 5.000 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.100 9.700 4.650 10.300 ;
    END
  END x
END nand2_0

MACRO mx4_5
  CLASS  CORE ;
  FOREIGN mx4_5 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 22.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 22.500 2.500 ;
    END
  END vss!
  PIN d0
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 16.550 7.100 17.350 7.850 ;
        RECT 16.750 5.950 17.900 6.550 ;
        RECT 16.250 7.200 17.350 7.850 ;
        RECT 16.750 5.950 17.350 7.850 ;
    END
  END d0
  PIN d1
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 19.700 5.850 20.300 7.850 ;
    END
  END d1
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 22.500 16.250 ;
    END
  END vdd!
  PIN d2
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.700 5.950 5.800 6.550 ;
        RECT 5.200 7.250 6.550 7.850 ;
        RECT 5.200 7.100 5.950 7.850 ;
        RECT 5.200 5.950 5.800 7.850 ;
    END
  END d2
  PIN sl0
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 14.100 5.950 16.100 6.550 ;
    END
  END sl0
  PIN d3
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.200 5.850 2.800 7.850 ;
    END
  END d3
  PIN sl1
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 20.950 7.150 21.550 9.150 ;
    END
  END sl1
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 10.050 8.250 10.750 10.400 ;
        RECT 10.050 9.600 13.950 10.400 ;
    END
  END x
  PIN sl2
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.300 5.950 8.300 6.550 ;
    END
  END sl2
  PIN sl3
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.950 7.150 1.550 9.150 ;
    END
  END sl3
  OBS 
      LAYER Metal1 ;
        RECT 0.500 9.700 7.950 10.300 ;
        RECT 8.800 5.850 13.600 6.450 ;
        RECT 3.900 7.350 4.500 9.050 ;
        RECT 8.800 5.850 9.400 9.050 ;
        RECT 2.150 8.450 9.400 9.050 ;
        RECT 11.700 6.950 12.350 7.550 ;
        RECT 11.700 6.950 12.300 9.050 ;
        RECT 18.000 7.350 18.600 9.050 ;
        RECT 11.700 8.450 20.350 9.050 ;
        RECT 14.550 9.700 22.000 10.300 ;
  END 
END mx4_5

MACRO mx4_4
  CLASS  CORE ;
  FOREIGN mx4_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 21.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 21.250 2.500 ;
    END
  END vss!
  PIN d0
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 17.250 5.950 19.250 6.550 ;
    END
  END d0
  PIN d1
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 15.000 7.200 17.000 7.800 ;
    END
  END d1
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 21.250 16.250 ;
    END
  END vdd!
  PIN d2
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.200 5.900 2.800 7.900 ;
    END
  END d2
  PIN sl0
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 18.700 8.450 20.700 9.050 ;
    END
  END sl0
  PIN d3
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.650 7.200 5.650 7.800 ;
    END
  END d3
  PIN sl1
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 12.500 7.200 14.500 7.800 ;
    END
  END sl1
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.350 9.700 11.750 10.300 ;
    END
  END x
  PIN sl2
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.350 8.450 2.350 9.050 ;
    END
  END sl2
  PIN sl3
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.400 7.200 8.400 7.800 ;
    END
  END sl3
  OBS 
      LAYER Metal1 ;
        RECT 0.450 9.700 7.850 10.300 ;
        RECT 3.250 4.800 13.150 5.400 ;
        RECT 8.900 4.800 9.500 9.050 ;
        RECT 5.550 8.450 9.500 9.050 ;
        RECT 13.750 4.850 17.850 5.450 ;
        RECT 13.750 4.850 14.350 6.500 ;
        RECT 11.400 5.900 14.350 6.500 ;
        RECT 11.400 5.900 12.000 9.050 ;
        RECT 11.400 8.450 15.550 9.050 ;
        RECT 13.250 9.700 20.650 10.300 ;
  END 
END mx4_4

MACRO mx4_3
  CLASS  CORE ;
  FOREIGN mx4_3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 21.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 21.250 2.500 ;
    END
  END vss!
  PIN d0
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.200 5.850 2.800 7.850 ;
    END
  END d0
  PIN d1
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.750 7.200 5.750 7.800 ;
    END
  END d1
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 21.250 16.250 ;
    END
  END vdd!
  PIN d2
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 18.450 5.850 19.050 7.850 ;
    END
  END d2
  PIN sl0
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.400 8.350 1.850 9.200 ;
    END
  END sl0
  PIN d3
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 15.100 7.200 17.100 7.800 ;
    END
  END d3
  PIN sl1
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.350 7.200 8.350 7.800 ;
    END
  END sl1
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.600 5.950 11.650 6.550 ;
    END
  END x
  PIN sl2
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 18.750 8.450 20.750 9.050 ;
    END
  END sl2
  PIN sl3
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 12.550 7.200 14.550 7.800 ;
    END
  END sl3
  OBS 
      LAYER Metal1 ;
        RECT 0.450 9.700 7.850 10.300 ;
        RECT 3.800 8.450 8.850 9.050 ;
        RECT 11.400 7.800 12.050 9.050 ;
        RECT 11.400 8.450 17.250 9.050 ;
        RECT 13.250 9.700 20.650 10.300 ;
  END 
END mx4_3

MACRO mx4_2
  CLASS  CORE ;
  FOREIGN mx4_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 21.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 21.250 2.500 ;
    END
  END vss!
  PIN d0
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.200 5.850 2.800 7.850 ;
    END
  END d0
  PIN d1
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.800 7.200 5.800 7.800 ;
    END
  END d1
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 21.250 16.250 ;
    END
  END vdd!
  PIN d2
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 18.450 5.850 19.050 7.850 ;
    END
  END d2
  PIN sl0
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.400 8.450 2.400 9.050 ;
    END
  END sl0
  PIN d3
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 15.250 7.200 17.250 7.800 ;
    END
  END d3
  PIN sl1
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.350 7.200 8.350 7.800 ;
    END
  END sl1
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.600 5.950 11.600 6.550 ;
    END
  END x
  PIN sl2
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 18.700 8.450 20.700 9.050 ;
    END
  END sl2
  PIN sl3
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 12.750 7.200 14.750 7.800 ;
    END
  END sl3
  OBS 
      LAYER Metal1 ;
        RECT 0.450 9.700 7.850 10.300 ;
        RECT 3.800 8.450 8.800 9.050 ;
        RECT 11.800 8.450 17.250 9.050 ;
        RECT 13.250 9.700 20.650 10.300 ;
  END 
END mx4_2

MACRO mx4_1
  CLASS  CORE ;
  FOREIGN mx4_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 17.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 17.500 2.500 ;
    END
  END vss!
  PIN d0
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 15.750 7.100 17.250 7.900 ;
    END
  END d0
  PIN d1
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 13.400 4.700 15.400 5.300 ;
    END
  END d1
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 17.500 16.250 ;
    END
  END vdd!
  PIN d2
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 7.100 1.750 7.900 ;
    END
  END d2
  PIN sl0
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.650 7.200 11.650 7.800 ;
    END
  END sl0
  PIN d3
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.600 4.700 3.600 5.300 ;
    END
  END d3
  PIN sl1
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 12.150 7.200 14.150 7.800 ;
    END
  END sl1
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.350 4.700 10.400 5.300 ;
    END
  END x
  PIN sl2
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.600 7.200 8.050 7.800 ;
    END
  END sl2
  PIN sl3
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.500 5.950 5.500 6.550 ;
    END
  END sl3
  OBS 
      LAYER Metal1 ;
        RECT 1.500 5.950 2.850 6.550 ;
        RECT 2.250 5.950 2.850 9.050 ;
        RECT 1.250 8.450 7.500 9.050 ;
        RECT 14.650 5.900 15.950 6.500 ;
        RECT 14.650 5.900 15.250 9.050 ;
        RECT 9.200 8.450 16.200 9.050 ;
  END 
END mx4_1

MACRO mux4_5
  CLASS  CORE ;
  FOREIGN mux4_5 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 28.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 28.750 2.500 ;
    END
  END vss!
  PIN d0
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 24.600 7.100 28.500 7.900 ;
    END
  END d0
  PIN d1
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 19.500 7.100 21.650 7.900 ;
    END
  END d1
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 28.750 16.250 ;
    END
  END vdd!
  PIN d2
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.450 5.950 3.900 6.550 ;
    END
  END d2
  PIN sl0
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.450 8.450 4.650 9.050 ;
    END
  END sl0
  PIN d3
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.100 7.100 9.100 7.900 ;
    END
  END d3
  PIN sl1
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.600 6.950 10.900 7.950 ;
    END
  END sl1
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 14.600 5.850 17.400 6.650 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 5.600 5.850 12.000 6.450 ;
        RECT 11.400 5.850 12.000 9.050 ;
        RECT 5.600 8.450 12.000 9.050 ;
        RECT 18.200 6.400 18.800 7.800 ;
        RECT 12.500 7.200 18.800 7.800 ;
        RECT 12.500 6.050 13.100 8.700 ;
        RECT 22.500 6.450 23.100 9.050 ;
        RECT 14.200 8.450 23.100 9.050 ;
        RECT 0.300 4.700 27.800 5.300 ;
        RECT 4.400 4.700 5.000 7.850 ;
        RECT 4.400 7.250 5.600 7.850 ;
        RECT 0.300 4.700 0.900 10.250 ;
        RECT 0.300 9.650 1.100 10.250 ;
  END 
END mux4_5

MACRO mux4_4
  CLASS  CORE ;
  FOREIGN mux4_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 28.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 28.750 2.500 ;
    END
  END vss!
  PIN d0
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 24.600 7.100 28.500 7.900 ;
    END
  END d0
  PIN d1
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 19.500 7.100 21.650 7.900 ;
    END
  END d1
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 28.750 16.250 ;
    END
  END vdd!
  PIN d2
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.450 5.950 3.900 6.550 ;
    END
  END d2
  PIN sl0
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.450 8.450 4.650 9.050 ;
    END
  END sl0
  PIN d3
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.100 7.100 9.100 7.900 ;
    END
  END d3
  PIN sl1
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.600 6.950 10.900 7.950 ;
    END
  END sl1
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 14.600 5.850 17.400 6.650 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 5.600 5.850 12.000 6.450 ;
        RECT 11.400 5.850 12.000 9.050 ;
        RECT 5.600 8.450 12.000 9.050 ;
        RECT 18.200 6.400 18.800 7.800 ;
        RECT 12.500 7.200 18.800 7.800 ;
        RECT 12.500 6.050 13.100 8.700 ;
        RECT 22.500 6.450 23.100 9.050 ;
        RECT 14.200 8.450 23.100 9.050 ;
        RECT 0.300 4.700 27.800 5.300 ;
        RECT 4.400 4.700 5.000 7.850 ;
        RECT 4.400 7.250 5.600 7.850 ;
        RECT 0.300 4.700 0.900 10.250 ;
        RECT 0.300 9.650 1.100 10.250 ;
  END 
END mux4_4

MACRO mux4_3
  CLASS  CORE ;
  FOREIGN mux4_3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 27.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 27.500 2.500 ;
    END
  END vss!
  PIN d0
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 23.750 7.200 25.750 7.800 ;
    END
  END d0
  PIN d1
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 18.750 7.200 20.850 7.800 ;
    END
  END d1
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 27.500 16.250 ;
    END
  END vdd!
  PIN d2
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.450 7.200 5.450 7.800 ;
    END
  END d2
  PIN sl0
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.300 8.450 2.300 9.050 ;
    END
  END sl0
  PIN d3
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.450 5.850 9.050 7.800 ;
        RECT 8.450 7.200 10.350 7.800 ;
    END
  END d3
  PIN sl1
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 10.950 7.050 11.550 9.050 ;
    END
  END sl1
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 15.050 5.950 18.250 6.550 ;
        RECT 16.650 8.450 18.250 9.050 ;
        RECT 17.650 5.950 18.250 9.050 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 11.950 5.800 13.150 6.400 ;
        RECT 6.750 6.450 7.350 10.300 ;
        RECT 12.550 5.800 13.150 10.300 ;
        RECT 6.750 9.700 13.150 10.300 ;
        RECT 13.650 7.150 17.050 7.750 ;
        RECT 13.650 6.050 14.250 8.700 ;
        RECT 3.300 4.700 18.950 5.300 ;
        RECT 21.750 6.450 22.350 10.300 ;
        RECT 15.350 9.700 22.350 10.300 ;
  END 
END mux4_3

MACRO mux4_2
  CLASS  CORE ;
  FOREIGN mux4_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 27.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 27.500 2.500 ;
    END
  END vss!
  PIN d0
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 23.750 7.200 25.750 7.800 ;
    END
  END d0
  PIN d1
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 18.750 7.200 20.850 7.800 ;
    END
  END d1
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 27.500 16.250 ;
    END
  END vdd!
  PIN d2
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.450 7.200 5.450 7.800 ;
    END
  END d2
  PIN sl0
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.300 8.450 2.300 9.050 ;
    END
  END sl0
  PIN d3
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.350 7.200 10.350 7.800 ;
    END
  END d3
  PIN sl1
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 10.850 6.450 11.650 7.900 ;
        RECT 10.850 7.100 12.050 7.900 ;
    END
  END sl1
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 15.050 5.950 18.150 6.550 ;
        RECT 16.650 8.300 18.150 8.900 ;
        RECT 17.550 5.950 18.150 8.900 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 3.350 5.050 10.800 5.650 ;
        RECT 11.950 5.050 13.150 5.650 ;
        RECT 6.700 6.450 7.400 10.000 ;
        RECT 12.550 5.050 13.150 10.000 ;
        RECT 6.700 9.400 13.150 10.000 ;
        RECT 13.650 7.200 17.050 7.800 ;
        RECT 13.650 6.450 14.250 9.100 ;
        RECT 21.750 6.450 22.350 10.000 ;
        RECT 15.350 9.400 22.350 10.000 ;
  END 
END mux4_2

MACRO mux4_1
  CLASS  CORE ;
  FOREIGN mux4_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 25.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 25.000 2.500 ;
    END
  END vss!
  PIN d0
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 22.400 8.450 24.400 9.050 ;
    END
  END d0
  PIN d1
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 17.050 7.200 19.150 7.800 ;
    END
  END d1
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 25.000 16.250 ;
    END
  END vdd!
  PIN d2
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.200 7.200 4.200 7.800 ;
    END
  END d2
  PIN sl0
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 8.450 2.250 9.050 ;
    END
  END sl0
  PIN d3
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.000 8.450 9.000 9.050 ;
    END
  END d3
  PIN sl1
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.600 5.950 10.600 6.550 ;
    END
  END sl1
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 13.350 5.950 16.550 6.550 ;
        RECT 14.950 8.700 16.550 9.300 ;
        RECT 15.950 5.950 16.550 9.300 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 5.050 6.450 5.650 10.400 ;
        RECT 5.050 9.800 10.850 10.400 ;
        RECT 11.950 7.200 15.350 7.800 ;
        RECT 11.950 6.450 12.550 9.100 ;
        RECT 20.050 6.450 20.650 10.400 ;
        RECT 13.650 9.800 20.650 10.400 ;
        RECT 21.150 5.950 22.350 6.550 ;
        RECT 21.150 5.950 21.750 10.400 ;
        RECT 21.150 9.800 22.350 10.400 ;
  END 
END mux4_1

MACRO mux2i_8
  CLASS  CORE ;
  FOREIGN mux2i_8 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 30.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 5.150 0.000 5.750 2.800 ;
        RECT 0.000 0.000 30.000 2.500 ;
    END
  END vss!
  PIN d0
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.350 5.950 6.450 6.550 ;
    END
  END d0
  PIN d1
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 22.000 5.950 24.250 6.550 ;
    END
  END d1
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 30.000 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 11.950 8.450 19.350 9.050 ;
    END
  END x
  PIN sl
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.950 4.700 1.550 5.550 ;
        RECT 8.450 5.950 17.200 6.550 ;
        RECT 8.450 4.700 9.050 6.550 ;
        RECT 0.950 4.700 9.050 5.300 ;
    END
  END sl
  OBS 
      LAYER Metal1 ;
        RECT 3.450 9.700 14.250 10.300 ;
        RECT 10.250 4.550 14.250 5.150 ;
        RECT 2.150 7.200 17.250 7.800 ;
        RECT 16.600 7.200 17.250 7.950 ;
        RECT 17.050 9.700 27.850 10.300 ;
        RECT 17.050 4.700 27.850 5.300 ;
  END 
END mux2i_8

MACRO mux2i_6
  CLASS  CORE ;
  FOREIGN mux2i_6 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 25.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 25.000 2.500 ;
    END
  END vss!
  PIN d0
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.550 5.950 3.150 7.900 ;
        RECT 1.400 7.100 3.150 7.900 ;
    END
  END d0
  PIN d1
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 18.850 5.950 21.200 6.550 ;
    END
  END d1
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 25.000 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.050 8.450 16.450 9.050 ;
    END
  END x
  PIN sl
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.400 4.700 2.000 6.550 ;
        RECT 12.250 5.900 14.150 6.550 ;
        RECT 9.700 5.650 12.850 6.250 ;
        RECT 9.850 5.650 10.450 6.600 ;
        RECT 5.950 5.950 10.450 6.550 ;
        RECT 5.950 4.700 6.550 6.550 ;
        RECT 1.400 4.700 6.550 5.300 ;
        RECT 1.400 4.700 2.100 5.400 ;
    END
  END sl
  OBS 
      LAYER Metal1 ;
        RECT 3.850 9.700 11.350 10.300 ;
        RECT 7.250 4.550 11.350 5.150 ;
        RECT 11.000 6.800 11.600 7.800 ;
        RECT 7.300 7.200 14.250 7.800 ;
        RECT 0.300 4.550 0.900 9.050 ;
        RECT 7.300 7.200 7.900 9.050 ;
        RECT 0.300 8.450 7.900 9.050 ;
        RECT 14.150 9.700 21.150 10.300 ;
        RECT 14.150 4.700 21.150 5.300 ;
  END 
END mux2i_6

MACRO mux2i_5
  CLASS  CORE ;
  FOREIGN mux2i_5 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 23.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 2.150 0.000 2.750 2.800 ;
        RECT 0.000 0.000 23.750 2.500 ;
    END
  END vss!
  PIN d0
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.550 7.200 3.550 7.800 ;
    END
  END d0
  PIN d1
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 18.350 5.950 20.700 6.550 ;
    END
  END d1
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 23.750 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.550 8.450 15.950 9.050 ;
    END
  END x
  PIN sl
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.850 5.950 14.000 6.550 ;
    END
  END sl
  OBS 
      LAYER Metal1 ;
        RECT 0.450 9.700 10.850 10.300 ;
        RECT 0.450 4.700 10.850 5.300 ;
        RECT 7.250 7.250 13.800 7.850 ;
        RECT 13.650 9.700 20.650 10.300 ;
        RECT 13.650 4.700 20.650 5.300 ;
  END 
END mux2i_5

MACRO mux2i_4
  CLASS  CORE ;
  FOREIGN mux2i_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 20.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 20.000 2.500 ;
    END
  END vss!
  PIN d0
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.550 5.950 3.350 7.900 ;
        RECT 2.100 7.100 3.350 7.900 ;
    END
  END d0
  PIN d1
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 16.650 5.950 18.650 6.550 ;
    END
  END d1
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 20.000 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 13.950 5.700 15.650 6.300 ;
        RECT 7.150 8.450 15.650 9.050 ;
        RECT 15.050 5.700 15.650 9.050 ;
    END
  END x
  PIN sl
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.400 4.700 2.000 6.550 ;
        RECT 10.950 5.800 12.250 6.400 ;
        RECT 5.950 5.650 11.550 6.250 ;
        RECT 5.950 4.700 6.650 6.250 ;
        RECT 1.400 4.700 6.650 5.300 ;
        RECT 1.400 4.700 2.100 5.400 ;
    END
  END sl
  OBS 
      LAYER Metal1 ;
        RECT 4.000 9.700 9.450 10.300 ;
        RECT 0.250 4.700 0.900 5.300 ;
        RECT 9.250 6.750 9.850 7.800 ;
        RECT 13.750 6.800 14.350 7.800 ;
        RECT 5.550 7.200 14.350 7.800 ;
        RECT 0.250 4.700 0.850 9.050 ;
        RECT 5.550 7.200 6.150 9.050 ;
        RECT 0.250 8.450 6.150 9.050 ;
        RECT 12.250 4.600 19.750 5.200 ;
        RECT 19.150 4.600 19.750 10.300 ;
        RECT 12.250 9.700 19.750 10.300 ;
  END 
END mux2i_4

MACRO mux2i_3
  CLASS  CORE ;
  FOREIGN mux2i_3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 15.000 2.500 ;
    END
  END vss!
  PIN d0
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.750 7.200 2.750 7.800 ;
    END
  END d0
  PIN d1
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 12.150 5.950 14.350 6.550 ;
    END
  END d1
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 15.000 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.400 7.200 10.400 7.800 ;
    END
  END x
  PIN sl
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.200 5.950 10.300 6.550 ;
    END
  END sl
  OBS 
      LAYER Metal1 ;
        RECT 2.200 8.450 7.500 9.050 ;
        RECT 2.200 4.700 7.500 5.300 ;
        RECT 10.300 4.650 14.300 5.250 ;
        RECT 10.900 4.650 11.500 9.050 ;
        RECT 10.300 8.450 14.300 9.050 ;
  END 
END mux2i_3

MACRO mux2i_2
  CLASS  CORE ;
  FOREIGN mux2i_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 12.500 2.500 ;
    END
  END vss!
  PIN d0
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.650 5.950 4.650 6.550 ;
    END
  END d0
  PIN d1
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.000 5.950 11.000 6.550 ;
    END
  END d1
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 9.650 13.450 10.250 16.250 ;
        RECT 0.000 13.750 12.500 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.300 8.450 7.400 9.050 ;
    END
  END x
  PIN sl
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 4.700 2.150 5.300 ;
        RECT 1.350 7.200 5.750 7.800 ;
        RECT 5.150 6.100 5.750 7.800 ;
        RECT 1.550 4.700 2.150 7.800 ;
    END
  END sl
  OBS 
      LAYER Metal1 ;
        RECT 0.250 6.050 1.000 6.650 ;
        RECT 0.250 6.050 0.850 9.150 ;
        RECT 0.250 8.550 1.050 9.150 ;
        RECT 6.250 4.700 6.850 7.800 ;
        RECT 7.950 8.450 11.950 9.050 ;
  END 
END mux2i_2

MACRO mux2i_1
  CLASS  CORE ;
  FOREIGN mux2i_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 10.000 2.500 ;
    END
  END vss!
  PIN d0
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.150 8.450 5.300 9.050 ;
    END
  END d0
  PIN d1
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.350 7.200 9.350 7.800 ;
    END
  END d1
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 10.000 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.550 9.700 7.900 10.300 ;
    END
  END x
  PIN sl
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.350 7.200 5.600 7.800 ;
    END
  END sl
  OBS 
      LAYER Metal1 ;
        RECT 0.250 5.950 0.950 6.550 ;
        RECT 0.250 5.950 0.850 9.450 ;
        RECT 0.250 8.800 1.050 9.450 ;
        RECT 5.550 5.950 6.700 6.550 ;
        RECT 6.100 5.950 6.700 9.100 ;
  END 
END mux2i_1

MACRO mux2_8
  CLASS  CORE ;
  FOREIGN mux2_8 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 15.000 2.500 ;
    END
  END vss!
  PIN d0
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.250 5.950 4.250 6.550 ;
    END
  END d0
  PIN d1
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.250 5.950 9.250 6.550 ;
    END
  END d1
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 15.000 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 10.500 7.200 14.600 7.800 ;
    END
  END x
  PIN sl
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.450 8.450 5.500 9.050 ;
    END
  END sl
  OBS 
      LAYER Metal1 ;
        RECT 4.900 6.600 5.500 7.800 ;
        RECT 0.350 7.150 5.500 7.800 ;
        RECT 0.350 5.950 0.950 10.300 ;
        RECT 0.350 9.700 1.050 10.300 ;
        RECT 5.450 5.500 6.600 6.100 ;
        RECT 6.000 8.400 13.500 9.100 ;
        RECT 6.000 5.500 6.600 10.300 ;
        RECT 5.450 9.700 6.600 10.300 ;
  END 
END mux2_8

MACRO mux2_6
  CLASS  CORE ;
  FOREIGN mux2_6 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 13.750 2.500 ;
    END
  END vss!
  PIN d0
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.150 5.950 4.150 6.550 ;
    END
  END d0
  PIN d1
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.500 5.950 9.500 6.550 ;
    END
  END d1
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 13.750 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 10.100 8.450 12.100 9.050 ;
    END
  END x
  PIN sl
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.350 8.450 3.350 9.050 ;
    END
  END sl
  OBS 
      LAYER Metal1 ;
        RECT 0.250 6.000 1.050 6.600 ;
        RECT 0.250 7.200 5.600 7.800 ;
        RECT 0.250 6.000 0.850 10.200 ;
        RECT 0.250 9.600 1.050 10.200 ;
        RECT 5.550 5.950 6.700 6.550 ;
        RECT 6.100 7.150 12.550 7.850 ;
        RECT 6.100 5.950 6.700 10.300 ;
        RECT 5.550 9.700 6.700 10.300 ;
  END 
END mux2_6

MACRO mux2_5
  CLASS  CORE ;
  FOREIGN mux2_5 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 13.750 2.500 ;
    END
  END vss!
  PIN d0
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.600 8.450 3.600 9.050 ;
    END
  END d0
  PIN d1
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.650 5.950 9.650 6.550 ;
    END
  END d1
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 2.150 13.550 2.750 16.250 ;
        RECT 0.000 13.750 13.750 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 10.100 8.450 12.100 9.050 ;
    END
  END x
  PIN sl
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.550 5.950 4.150 6.550 ;
    END
  END sl
  OBS 
      LAYER Metal1 ;
        RECT 0.450 7.200 5.600 7.800 ;
        RECT 0.450 4.850 1.050 9.150 ;
        RECT 5.550 5.950 6.700 6.550 ;
        RECT 6.100 7.150 12.550 7.850 ;
        RECT 6.100 5.950 6.700 9.050 ;
        RECT 5.550 8.450 6.700 9.050 ;
  END 
END mux2_5

MACRO mux2_4
  CLASS  CORE ;
  FOREIGN mux2_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 12.500 2.500 ;
    END
  END vss!
  PIN d0
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.150 5.950 4.150 6.550 ;
    END
  END d0
  PIN d1
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.100 5.950 9.100 6.550 ;
    END
  END d1
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 12.500 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.850 8.500 12.150 9.100 ;
    END
  END x
  PIN sl
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.450 8.450 3.450 9.050 ;
    END
  END sl
  OBS 
      LAYER Metal1 ;
        RECT 4.600 6.950 5.200 7.800 ;
        RECT 0.350 7.200 5.200 7.800 ;
        RECT 0.350 5.850 0.950 10.300 ;
        RECT 0.350 9.700 1.050 10.300 ;
        RECT 5.150 5.850 6.300 6.450 ;
        RECT 5.700 7.150 9.200 7.850 ;
        RECT 8.600 7.150 9.200 7.900 ;
        RECT 5.700 5.850 6.300 10.300 ;
        RECT 5.150 9.700 6.300 10.300 ;
  END 
END mux2_4

MACRO mux2_3
  CLASS  CORE ;
  FOREIGN mux2_3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 12.500 2.500 ;
    END
  END vss!
  PIN d0
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.500 8.450 3.500 9.050 ;
    END
  END d0
  PIN d1
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.100 5.950 9.100 6.550 ;
    END
  END d1
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 1.750 13.550 2.350 16.250 ;
        RECT 0.000 13.750 12.500 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.850 8.450 12.000 9.050 ;
    END
  END x
  PIN sl
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.550 5.950 4.150 6.550 ;
    END
  END sl
  OBS 
      LAYER Metal1 ;
        RECT 0.350 7.200 5.200 7.800 ;
        RECT 0.350 4.700 0.950 9.150 ;
        RECT 5.150 5.950 6.300 6.550 ;
        RECT 5.700 7.150 9.600 7.850 ;
        RECT 5.700 5.950 6.300 9.050 ;
        RECT 5.150 8.450 6.300 9.050 ;
  END 
END mux2_3

MACRO mux2_2
  CLASS  CORE ;
  FOREIGN mux2_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 11.250 2.500 ;
    END
  END vss!
  PIN d0
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.200 7.200 4.200 7.800 ;
    END
  END d0
  PIN d1
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.000 5.950 9.000 6.550 ;
    END
  END d1
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 11.250 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.000 7.200 11.000 7.800 ;
    END
  END x
  PIN sl
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 8.450 2.250 9.050 ;
    END
  END sl
  OBS 
      LAYER Metal1 ;
        RECT 5.000 6.450 5.700 9.100 ;
        RECT 5.000 8.400 9.700 9.100 ;
  END 
END mux2_2

MACRO mux2_1
  CLASS  CORE ;
  FOREIGN mux2_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 11.250 2.500 ;
    END
  END vss!
  PIN d0
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.200 7.200 4.200 7.800 ;
    END
  END d0
  PIN d1
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.000 5.950 9.000 6.550 ;
    END
  END d1
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 11.250 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.000 7.200 11.000 7.800 ;
    END
  END x
  PIN sl
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 8.450 2.250 9.050 ;
    END
  END sl
  OBS 
      LAYER Metal1 ;
        RECT 4.950 6.450 5.650 9.100 ;
        RECT 4.950 8.400 9.450 9.100 ;
  END 
END mux2_1

MACRO latpr_8
  CLASS  CORE ;
  FOREIGN latpr_8 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 23.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 18.150 9.700 20.150 10.300 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 23.750 2.500 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.900 8.450 2.900 9.050 ;
    END
  END d
  PIN gb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 21.300 5.950 23.450 6.550 ;
    END
  END gb
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 3.050 13.450 3.650 16.250 ;
        RECT 0.000 13.750 23.750 16.250 ;
        RECT 13.900 13.450 14.500 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 14.600 9.700 16.600 10.300 ;
    END
  END qb
  PIN rb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.950 5.850 1.550 7.850 ;
    END
  END rb
  OBS 
      LAYER Metal1 ;
        RECT 1.350 9.700 5.350 10.300 ;
        RECT 5.950 7.350 11.500 7.950 ;
        RECT 8.800 6.100 12.800 6.700 ;
        RECT 5.000 4.650 5.600 5.600 ;
        RECT 3.650 5.000 5.600 5.600 ;
        RECT 13.300 6.100 18.300 6.700 ;
        RECT 3.650 5.000 4.250 9.150 ;
        RECT 13.300 6.100 13.900 9.150 ;
        RECT 3.650 8.550 13.900 9.150 ;
        RECT 7.000 8.550 7.650 9.200 ;
        RECT 9.150 4.750 9.750 5.600 ;
        RECT 7.250 5.000 20.350 5.600 ;
        RECT 7.250 5.000 7.850 6.850 ;
        RECT 4.800 6.250 7.850 6.850 ;
        RECT 19.750 5.000 20.350 7.800 ;
        RECT 19.750 7.200 23.000 7.800 ;
  END 
END latpr_8

MACRO latpr_4
  CLASS  CORE ;
  FOREIGN latpr_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 20.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 10.750 8.450 12.900 9.050 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 8.200 0.000 8.800 2.800 ;
        RECT 0.000 0.000 20.000 2.500 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.750 8.450 2.900 9.050 ;
    END
  END d
  PIN gb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 17.100 5.950 19.250 6.550 ;
    END
  END gb
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 20.000 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 14.500 8.450 16.750 9.050 ;
    END
  END qb
  PIN rb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.100 4.700 8.050 5.300 ;
    END
  END rb
  OBS 
      LAYER Metal1 ;
        RECT 5.050 8.600 9.200 9.200 ;
        RECT 9.850 4.700 13.900 5.300 ;
        RECT 5.450 5.800 6.050 6.550 ;
        RECT 5.450 5.950 16.500 6.550 ;
        RECT 4.050 6.750 4.700 7.800 ;
        RECT 4.050 7.200 19.650 7.800 ;
  END 
END latpr_4

MACRO latpr_2
  CLASS  CORE ;
  FOREIGN latpr_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 16.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.750 5.950 11.750 6.550 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 9.100 0.000 9.700 2.700 ;
        RECT 0.000 0.000 16.250 2.500 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.300 7.200 3.300 7.800 ;
    END
  END d
  PIN gb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 14.000 8.450 16.000 9.050 ;
    END
  END gb
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 3.650 13.550 4.250 16.250 ;
        RECT 0.000 13.750 16.250 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.550 5.950 8.550 6.550 ;
    END
  END qb
  PIN rb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 3.450 8.200 4.050 ;
    END
  END rb
  OBS 
      LAYER Metal1 ;
        RECT 4.250 6.050 4.850 9.050 ;
        RECT 4.250 8.450 13.500 9.050 ;
        RECT 5.750 7.250 14.800 7.850 ;
  END 
END latpr_2

MACRO latpr_1
  CLASS  CORE ;
  FOREIGN latpr_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.000 5.950 11.000 6.550 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 8.450 0.000 9.050 2.700 ;
        RECT 0.000 0.000 15.000 2.500 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.300 7.200 3.300 7.800 ;
    END
  END d
  PIN gb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 12.750 9.700 14.750 10.300 ;
    END
  END gb
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 1.250 13.550 1.850 16.250 ;
        RECT 0.000 13.750 15.000 16.250 ;
        RECT 8.150 13.450 8.750 16.250 ;
        RECT 3.050 13.550 3.650 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.000 5.950 8.000 6.550 ;
    END
  END qb
  PIN rb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 3.450 7.750 4.050 ;
    END
  END rb
  OBS 
      LAYER Metal1 ;
        RECT 4.050 6.150 4.850 6.750 ;
        RECT 4.050 6.150 4.650 9.050 ;
        RECT 4.050 8.450 12.250 9.050 ;
        RECT 5.200 7.250 13.850 7.850 ;
  END 
END latpr_1

MACRO latp_8
  CLASS  CORE ;
  FOREIGN latp_8 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 21.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 15.800 9.700 17.800 10.300 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.700 0.000 1.300 2.800 ;
        RECT 0.000 0.000 21.250 2.500 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.300 8.450 2.300 9.050 ;
    END
  END d
  PIN gb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 18.750 5.950 19.350 7.800 ;
        RECT 8.550 7.200 20.800 7.800 ;
        RECT 18.750 7.100 19.600 7.800 ;
    END
  END gb
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 11.550 13.450 12.150 16.250 ;
        RECT 0.000 13.750 21.250 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 12.250 9.700 14.250 10.300 ;
    END
  END qb
  OBS 
      LAYER Metal1 ;
        RECT 0.450 9.700 4.450 10.300 ;
        RECT 3.100 5.500 4.700 6.100 ;
        RECT 7.450 5.950 15.950 6.550 ;
        RECT 3.100 5.500 3.700 9.150 ;
        RECT 7.450 5.950 8.050 9.150 ;
        RECT 3.100 8.550 8.050 9.150 ;
        RECT 5.300 4.750 20.650 5.350 ;
        RECT 5.300 4.750 5.900 7.300 ;
        RECT 4.200 6.600 5.900 7.300 ;
        RECT 4.200 6.700 6.950 7.300 ;
  END 
END latp_8

MACRO latp_4
  CLASS  CORE ;
  FOREIGN latp_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 17.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.600 8.450 9.600 9.050 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 5.650 0.000 6.250 2.800 ;
        RECT 0.000 0.000 17.500 2.500 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.300 4.700 3.050 5.300 ;
    END
  END d
  PIN gb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 15.150 5.950 17.250 6.550 ;
    END
  END gb
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 5.650 13.450 6.250 16.250 ;
        RECT 0.000 13.750 17.500 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 11.200 8.450 13.200 9.050 ;
    END
  END qb
  OBS 
      LAYER Metal1 ;
        RECT 7.350 4.700 11.350 5.300 ;
        RECT 4.700 5.950 13.950 6.550 ;
        RECT 3.350 6.650 3.950 7.800 ;
        RECT 3.350 7.200 17.050 7.800 ;
  END 
END latp_4

MACRO latp_2
  CLASS  CORE ;
  FOREIGN latp_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.750 5.950 9.750 6.550 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 6.850 0.000 7.450 2.800 ;
        RECT 0.000 0.000 13.750 2.500 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 7.200 2.250 7.800 ;
    END
  END d
  PIN gb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 11.500 9.700 13.500 10.300 ;
    END
  END gb
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 6.950 13.450 7.550 16.250 ;
        RECT 0.000 13.750 13.750 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.750 5.950 6.750 6.550 ;
    END
  END qb
  OBS 
      LAYER Metal1 ;
        RECT 2.950 6.150 3.900 6.750 ;
        RECT 2.950 6.150 3.550 9.050 ;
        RECT 2.950 8.450 11.000 9.050 ;
        RECT 10.750 7.250 12.550 7.850 ;
        RECT 4.050 7.300 11.350 7.900 ;
  END 
END latp_2

MACRO latp_1
  CLASS  CORE ;
  FOREIGN latp_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.500 5.950 9.500 6.550 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 6.850 0.000 7.450 2.800 ;
        RECT 0.000 0.000 13.750 2.500 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 7.200 2.250 7.800 ;
    END
  END d
  PIN gb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 11.500 9.700 13.500 10.300 ;
    END
  END gb
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 13.750 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.750 5.950 6.750 6.550 ;
    END
  END qb
  OBS 
      LAYER Metal1 ;
        RECT 3.000 6.150 3.900 6.750 ;
        RECT 3.000 6.150 3.600 9.050 ;
        RECT 3.000 8.450 11.000 9.050 ;
        RECT 10.750 7.250 12.550 7.850 ;
        RECT 4.100 7.300 11.350 7.900 ;
  END 
END latp_1

MACRO latnr_8
  CLASS  CORE ;
  FOREIGN latnr_8 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 23.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 18.000 9.700 20.000 10.300 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 23.750 2.500 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.900 8.450 2.900 9.050 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 3.050 13.450 3.650 16.250 ;
        RECT 0.000 13.750 23.750 16.250 ;
        RECT 13.750 13.450 14.350 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 14.450 9.700 16.450 10.300 ;
    END
  END qb
  PIN g
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 20.950 5.950 23.200 6.550 ;
    END
  END g
  PIN rb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.950 5.850 1.550 7.850 ;
    END
  END rb
  OBS 
      LAYER Metal1 ;
        RECT 1.350 9.700 5.350 10.300 ;
        RECT 4.650 6.500 5.250 7.950 ;
        RECT 6.850 6.850 7.450 7.950 ;
        RECT 4.650 7.350 11.150 7.950 ;
        RECT 7.950 5.750 8.550 6.500 ;
        RECT 7.950 5.900 12.650 6.500 ;
        RECT 3.500 4.600 5.600 5.200 ;
        RECT 13.350 6.100 18.150 6.700 ;
        RECT 3.500 4.600 4.100 9.150 ;
        RECT 13.350 6.100 13.950 9.150 ;
        RECT 3.500 8.550 13.950 9.150 ;
        RECT 6.100 4.600 9.850 5.200 ;
        RECT 6.100 4.600 6.700 5.350 ;
        RECT 9.250 4.750 20.200 5.350 ;
        RECT 19.600 4.750 20.200 7.800 ;
        RECT 19.600 7.200 22.850 7.800 ;
  END 
END latnr_8

MACRO latnr_4
  CLASS  CORE ;
  FOREIGN latnr_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 20.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 10.100 8.450 12.100 9.050 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 8.150 0.000 8.750 2.800 ;
        RECT 0.000 0.000 20.000 2.500 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.400 8.450 2.400 9.050 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 20.000 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 13.700 8.450 15.700 9.050 ;
    END
  END qb
  PIN g
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 17.650 7.200 19.750 7.800 ;
    END
  END g
  PIN rb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.100 4.700 7.950 5.300 ;
    END
  END rb
  OBS 
      LAYER Metal1 ;
        RECT 2.950 5.900 3.550 9.050 ;
        RECT 5.450 8.450 9.050 9.200 ;
        RECT 9.850 4.700 13.850 5.300 ;
        RECT 4.150 6.600 4.750 7.800 ;
        RECT 4.150 7.200 16.450 7.800 ;
        RECT 5.450 5.950 19.550 6.550 ;
  END 
END latnr_4

MACRO latnr_2
  CLASS  CORE ;
  FOREIGN latnr_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 16.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.800 5.950 11.800 6.550 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 8.900 0.000 9.500 2.700 ;
        RECT 0.000 0.000 16.250 2.500 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.300 7.200 3.300 7.800 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 3.650 13.550 4.250 16.250 ;
        RECT 0.000 13.750 16.250 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.550 5.950 8.550 6.550 ;
    END
  END qb
  PIN g
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 13.950 5.950 15.950 6.550 ;
    END
  END g
  PIN rb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 3.450 8.200 4.050 ;
    END
  END rb
  OBS 
      LAYER Metal1 ;
        RECT 5.750 7.250 13.300 7.850 ;
        RECT 4.250 6.050 4.850 9.050 ;
        RECT 4.250 8.450 14.600 9.050 ;
  END 
END latnr_2

MACRO latnr_1
  CLASS  CORE ;
  FOREIGN latnr_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.000 5.950 11.000 6.550 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 8.450 0.000 9.050 2.700 ;
        RECT 0.000 0.000 15.000 2.500 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.300 7.200 3.300 7.800 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 1.250 13.550 1.850 16.250 ;
        RECT 0.000 13.750 15.000 16.250 ;
        RECT 8.150 13.450 8.750 16.250 ;
        RECT 3.050 13.550 3.650 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.000 5.950 8.000 6.550 ;
    END
  END qb
  PIN g
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 12.700 9.700 14.700 10.300 ;
    END
  END g
  PIN rb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 3.450 7.750 4.050 ;
    END
  END rb
  OBS 
      LAYER Metal1 ;
        RECT 5.200 7.250 12.250 7.850 ;
        RECT 4.050 6.150 4.850 6.750 ;
        RECT 4.050 6.150 4.650 9.050 ;
        RECT 4.050 8.450 13.350 9.050 ;
  END 
END latnr_1

MACRO latn_8
  CLASS  CORE ;
  FOREIGN latn_8 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 21.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 15.800 9.700 17.800 10.300 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.700 0.000 1.300 2.800 ;
        RECT 0.000 0.000 21.250 2.500 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 8.450 2.250 9.050 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 11.550 13.450 12.150 16.250 ;
        RECT 0.000 13.750 21.250 16.250 ;
        RECT 18.350 13.450 18.950 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 12.250 9.700 14.250 10.300 ;
    END
  END qb
  PIN g
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 18.650 5.950 20.650 6.550 ;
    END
  END g
  OBS 
      LAYER Metal1 ;
        RECT 2.400 6.300 3.350 6.900 ;
        RECT 2.750 6.300 3.350 10.300 ;
        RECT 0.450 9.700 4.450 10.300 ;
        RECT 4.950 6.700 5.550 7.450 ;
        RECT 4.950 6.850 7.600 7.450 ;
        RECT 3.850 5.600 4.700 6.200 ;
        RECT 10.950 6.100 15.950 6.700 ;
        RECT 3.850 5.600 4.450 9.150 ;
        RECT 10.950 6.100 11.550 9.150 ;
        RECT 3.850 8.550 11.550 9.150 ;
        RECT 6.300 5.000 18.000 5.600 ;
        RECT 6.300 5.000 6.900 6.200 ;
        RECT 17.400 5.000 18.000 7.800 ;
        RECT 17.400 7.200 20.650 7.800 ;
  END 
END latn_8

MACRO latn_4
  CLASS  CORE ;
  FOREIGN latn_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 17.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.600 8.450 9.600 9.050 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 5.650 0.000 6.250 2.800 ;
        RECT 0.000 0.000 17.500 2.500 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.300 4.700 3.050 5.300 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 5.650 13.450 6.250 16.250 ;
        RECT 0.000 13.750 17.500 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 11.200 8.450 13.200 9.050 ;
    END
  END qb
  PIN g
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 15.150 7.200 17.250 7.800 ;
    END
  END g
  OBS 
      LAYER Metal1 ;
        RECT 7.350 4.700 11.350 5.300 ;
        RECT 3.200 6.950 3.800 7.800 ;
        RECT 3.200 7.200 13.950 7.800 ;
        RECT 6.050 5.950 17.050 6.550 ;
  END 
END latn_4

MACRO latn_2
  CLASS  CORE ;
  FOREIGN latn_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.750 5.950 9.750 6.550 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 6.850 0.000 7.450 2.800 ;
        RECT 0.000 0.000 13.750 2.500 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 7.200 2.250 7.800 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 6.950 13.450 7.550 16.250 ;
        RECT 0.000 13.750 13.750 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.750 5.950 6.750 6.550 ;
    END
  END qb
  PIN g
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 11.400 9.700 13.400 10.300 ;
    END
  END g
  OBS 
      LAYER Metal1 ;
        RECT 4.050 7.300 11.000 7.900 ;
        RECT 2.950 6.150 3.900 6.750 ;
        RECT 2.950 6.150 3.550 9.050 ;
        RECT 2.950 8.450 12.100 9.050 ;
  END 
END latn_2

MACRO latn_1
  CLASS  CORE ;
  FOREIGN latn_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.750 5.950 9.750 6.550 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 6.850 0.000 7.450 2.800 ;
        RECT 0.000 0.000 13.750 2.500 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 7.200 2.250 7.800 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 13.750 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.750 5.950 6.750 6.550 ;
    END
  END qb
  PIN g
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 11.400 9.700 13.400 10.300 ;
    END
  END g
  OBS 
      LAYER Metal1 ;
        RECT 4.100 7.300 11.000 7.900 ;
        RECT 3.000 6.150 3.900 6.750 ;
        RECT 3.000 6.150 3.600 9.050 ;
        RECT 3.000 8.450 12.100 9.050 ;
  END 
END latn_1

MACRO inv_8
  CLASS  CORE ;
  FOREIGN inv_8 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.850 8.450 6.200 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 7.500 2.500 ;
    END
  END vss!
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 7.500 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.100 10.950 6.650 11.550 ;
    END
  END x
END inv_8

MACRO inv_7
  CLASS  CORE ;
  FOREIGN inv_7 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.850 8.450 5.600 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 7.500 2.500 ;
    END
  END vss!
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 7.500 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.100 10.950 6.650 11.550 ;
    END
  END x
END inv_7

MACRO inv_6
  CLASS  CORE ;
  FOREIGN inv_6 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.850 8.450 5.600 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 7.500 2.500 ;
    END
  END vss!
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 7.500 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.100 10.950 6.650 11.550 ;
    END
  END x
END inv_6

MACRO inv_5
  CLASS  CORE ;
  FOREIGN inv_5 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.800 8.450 4.100 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 5.000 2.500 ;
    END
  END vss!
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 5.000 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.250 5.950 3.250 6.550 ;
    END
  END x
END inv_5

MACRO inv_4
  CLASS  CORE ;
  FOREIGN inv_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.850 8.450 4.150 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 5.000 2.500 ;
    END
  END vss!
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 5.000 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.200 5.950 4.200 6.550 ;
    END
  END x
END inv_4

MACRO inv_3
  CLASS  CORE ;
  FOREIGN inv_3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.850 8.450 4.150 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 5.000 2.500 ;
    END
  END vss!
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 5.000 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.200 5.950 4.200 6.550 ;
    END
  END x
END inv_3

MACRO inv_2
  CLASS  CORE ;
  FOREIGN inv_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 8.450 2.250 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 3.750 2.500 ;
    END
  END vss!
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 3.750 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.500 5.950 3.500 6.550 ;
    END
  END x
END inv_2

MACRO inv_16
  CLASS  CORE ;
  FOREIGN inv_16 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.850 5.950 8.500 6.550 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 10.000 2.500 ;
    END
  END vss!
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 10.000 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.100 9.700 6.150 10.300 ;
    END
  END x
END inv_16

MACRO inv_14
  CLASS  CORE ;
  FOREIGN inv_14 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.850 7.200 8.450 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 10.000 2.500 ;
    END
  END vss!
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 10.000 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.150 9.700 6.150 10.300 ;
    END
  END x
END inv_14

MACRO inv_12
  CLASS  CORE ;
  FOREIGN inv_12 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.950 5.950 7.950 6.550 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 8.750 2.500 ;
    END
  END vss!
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 8.750 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.200 10.950 6.350 11.550 ;
    END
  END x
END inv_12

MACRO inv_10
  CLASS  CORE ;
  FOREIGN inv_10 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.950 7.200 6.450 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 8.750 2.500 ;
    END
  END vss!
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 8.750 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.200 10.950 6.350 11.550 ;
    END
  END x
END inv_10

MACRO inv_1
  CLASS  CORE ;
  FOREIGN inv_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 8.450 2.250 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 3.750 2.500 ;
    END
  END vss!
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 3.750 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.500 5.950 3.500 6.550 ;
    END
  END x
END inv_1

MACRO inv_0
  CLASS  CORE ;
  FOREIGN inv_0 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 8.450 2.250 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 3.750 2.500 ;
    END
  END vss!
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 3.750 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.500 5.950 3.500 6.550 ;
    END
  END x
END inv_0

MACRO exor3_5
  CLASS  CORE ;
  FOREIGN exor3_5 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 21.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.600 7.200 2.600 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 2.150 0.000 2.750 2.800 ;
        RECT 0.000 0.000 21.250 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.850 5.950 3.850 6.550 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.050 5.950 10.150 6.550 ;
    END
  END c
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 2.100 13.500 2.800 16.250 ;
        RECT 0.000 13.750 21.250 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 17.150 8.450 19.150 9.050 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 0.450 4.700 4.950 5.300 ;
        RECT 4.350 7.200 5.550 7.800 ;
        RECT 4.350 4.700 4.950 9.050 ;
        RECT 0.450 8.450 4.950 9.050 ;
        RECT 8.550 8.450 9.150 10.150 ;
        RECT 3.850 9.550 9.150 10.150 ;
        RECT 5.550 5.950 6.700 6.550 ;
        RECT 6.100 7.200 11.250 7.800 ;
        RECT 6.100 5.950 6.700 9.050 ;
        RECT 5.550 8.450 6.700 9.050 ;
        RECT 10.650 4.800 11.250 10.150 ;
        RECT 15.350 8.500 15.950 10.150 ;
        RECT 10.650 9.550 15.950 10.150 ;
        RECT 12.350 5.950 13.500 6.550 ;
        RECT 12.900 7.200 19.350 7.800 ;
        RECT 12.900 5.950 13.500 9.050 ;
        RECT 12.350 8.450 13.500 9.050 ;
  END 
END exor3_5

MACRO exor3_4
  CLASS  CORE ;
  FOREIGN exor3_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 20.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.750 7.200 2.750 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 2.150 0.000 2.750 2.800 ;
        RECT 0.000 0.000 20.000 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.150 5.950 3.150 6.550 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.400 5.950 10.400 6.550 ;
    END
  END c
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 2.100 13.500 2.800 16.250 ;
        RECT 0.000 13.750 20.000 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 17.200 8.450 19.250 9.050 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 0.450 4.700 4.950 5.300 ;
        RECT 4.350 7.200 5.550 7.800 ;
        RECT 4.350 4.700 4.950 9.050 ;
        RECT 0.450 8.450 4.950 9.050 ;
        RECT 8.550 8.450 9.150 10.150 ;
        RECT 3.850 9.550 9.150 10.150 ;
        RECT 10.650 4.700 11.500 5.300 ;
        RECT 5.550 5.950 6.700 6.550 ;
        RECT 10.900 4.700 11.500 7.800 ;
        RECT 6.100 7.200 11.500 7.800 ;
        RECT 6.100 5.950 6.700 9.050 ;
        RECT 5.550 8.450 6.700 9.050 ;
        RECT 10.650 7.200 11.250 10.150 ;
        RECT 15.350 8.000 15.950 10.150 ;
        RECT 10.650 9.550 15.950 10.150 ;
        RECT 12.350 6.900 19.150 7.500 ;
        RECT 12.350 5.950 12.950 9.050 ;
  END 
END exor3_4

MACRO exor3_3
  CLASS  CORE ;
  FOREIGN exor3_3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 18.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.850 7.200 2.850 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 2.150 0.000 2.750 2.800 ;
        RECT 0.000 0.000 18.750 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.150 5.950 3.150 6.550 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.400 5.950 10.400 6.550 ;
    END
  END c
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 2.100 13.500 2.800 16.250 ;
        RECT 0.000 13.750 18.750 16.250 ;
        RECT 15.850 13.100 16.450 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 17.650 4.700 18.400 5.300 ;
        RECT 17.200 8.450 18.400 9.050 ;
        RECT 17.800 4.700 18.400 9.050 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 0.450 4.700 4.950 5.300 ;
        RECT 4.350 7.200 5.550 7.800 ;
        RECT 4.350 4.700 4.950 9.050 ;
        RECT 0.450 8.450 4.950 9.050 ;
        RECT 8.550 8.450 9.150 10.150 ;
        RECT 3.850 9.550 9.150 10.150 ;
        RECT 10.650 4.700 11.500 5.300 ;
        RECT 5.550 5.950 6.700 6.550 ;
        RECT 10.900 5.950 15.950 6.550 ;
        RECT 10.900 4.700 11.500 7.800 ;
        RECT 6.100 7.200 11.500 7.800 ;
        RECT 6.100 5.950 6.700 9.050 ;
        RECT 5.550 8.450 6.700 9.050 ;
        RECT 10.650 7.200 11.250 10.150 ;
        RECT 12.350 4.700 17.050 5.300 ;
        RECT 16.450 5.950 17.300 6.550 ;
        RECT 16.450 4.700 17.050 7.800 ;
        RECT 12.350 7.200 17.050 7.800 ;
  END 
END exor3_3

MACRO exor3_2
  CLASS  CORE ;
  FOREIGN exor3_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 17.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.350 8.450 2.350 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 1.050 0.000 1.650 2.800 ;
        RECT 0.000 0.000 17.500 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.450 7.200 4.100 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.350 5.800 9.250 7.500 ;
    END
  END c
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 1.000 13.550 1.700 16.250 ;
        RECT 0.000 13.750 17.500 16.250 ;
        RECT 7.850 13.450 8.450 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 16.350 7.300 17.000 9.050 ;
        RECT 15.800 8.450 17.200 9.050 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 2.750 4.700 7.850 5.300 ;
        RECT 7.250 4.700 7.850 6.400 ;
        RECT 9.550 4.700 14.850 5.300 ;
        RECT 4.450 5.950 5.600 6.550 ;
        RECT 14.250 4.700 14.850 6.600 ;
        RECT 5.000 5.950 5.600 9.050 ;
        RECT 10.150 4.700 10.750 9.050 ;
        RECT 4.450 8.450 10.750 9.050 ;
        RECT 11.250 6.700 11.850 9.050 ;
        RECT 11.250 8.400 15.300 9.050 ;
  END 
END exor3_2

MACRO exor3_1
  CLASS  CORE ;
  FOREIGN exor3_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 17.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.350 8.450 2.350 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 1.000 0.000 1.600 2.800 ;
        RECT 0.000 0.000 17.500 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.800 5.950 2.800 6.550 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.500 5.950 9.500 6.550 ;
    END
  END c
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.950 13.550 1.650 16.250 ;
        RECT 0.000 13.750 17.500 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 15.950 7.400 16.550 9.050 ;
        RECT 15.950 8.450 16.900 9.050 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 2.700 4.700 6.800 5.300 ;
        RECT 6.200 4.700 6.800 7.800 ;
        RECT 6.200 7.200 8.000 7.800 ;
        RECT 9.500 4.700 14.800 5.300 ;
        RECT 14.200 4.700 14.800 6.700 ;
        RECT 4.400 5.950 5.000 9.050 ;
        RECT 10.000 4.700 10.600 9.050 ;
        RECT 4.400 8.450 10.600 9.050 ;
        RECT 11.200 8.100 15.200 8.700 ;
        RECT 11.200 5.950 11.800 9.050 ;
  END 
END exor3_1

MACRO exor2_8
  CLASS  CORE ;
  FOREIGN exor2_8 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 30.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.150 8.450 3.150 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 2.100 0.000 2.800 2.700 ;
        RECT 0.000 0.000 30.000 2.500 ;
        RECT 19.100 0.000 19.800 2.750 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.700 5.950 24.350 6.550 ;
    END
  END b
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 2.100 13.550 2.800 16.250 ;
        RECT 0.000 13.750 30.000 16.250 ;
        RECT 25.900 13.500 26.600 16.250 ;
        RECT 19.100 13.500 19.800 16.250 ;
        RECT 5.500 13.550 6.200 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.950 9.700 16.350 10.300 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 3.800 4.750 14.650 5.350 ;
        RECT 17.450 7.050 21.450 7.650 ;
        RECT 7.250 7.200 18.050 7.800 ;
        RECT 20.850 7.200 28.300 7.800 ;
        RECT 3.850 8.450 29.550 9.050 ;
  END 
END exor2_8

MACRO exor2_6
  CLASS  CORE ;
  FOREIGN exor2_6 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 23.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.150 8.450 3.150 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 2.100 0.000 2.800 2.700 ;
        RECT 0.000 0.000 23.750 2.500 ;
        RECT 20.800 0.000 21.500 2.750 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.700 5.950 9.650 6.550 ;
        RECT 12.200 5.950 16.600 6.550 ;
        RECT 9.050 5.750 12.800 6.350 ;
    END
  END b
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 2.100 13.550 2.800 16.250 ;
        RECT 0.000 13.750 23.750 16.250 ;
        RECT 19.100 13.500 19.800 16.250 ;
        RECT 15.700 13.500 16.400 16.250 ;
        RECT 5.500 13.550 6.200 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.950 9.700 12.950 10.300 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 3.850 8.450 18.050 9.050 ;
        RECT 10.650 6.850 11.250 7.800 ;
        RECT 7.250 7.200 21.450 7.800 ;
  END 
END exor2_6

MACRO exor2_5
  CLASS  CORE ;
  FOREIGN exor2_5 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 22.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.150 5.950 3.150 6.550 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 22.500 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.150 5.950 17.300 6.550 ;
    END
  END b
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 2.100 13.550 2.800 16.250 ;
        RECT 0.000 13.750 22.500 16.250 ;
        RECT 19.100 13.500 19.800 16.250 ;
        RECT 15.700 13.500 16.400 16.250 ;
        RECT 5.500 13.550 6.200 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.950 4.700 12.950 5.300 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 3.850 10.950 18.050 11.550 ;
        RECT 7.250 8.000 21.450 8.600 ;
  END 
END exor2_5

MACRO exor2_4
  CLASS  CORE ;
  FOREIGN exor2_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 18.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.200 6.950 2.800 7.800 ;
        RECT 0.950 7.200 2.800 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 2.350 0.000 3.050 2.700 ;
        RECT 0.000 0.000 18.750 2.500 ;
        RECT 15.950 0.000 16.650 2.800 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.700 5.950 4.700 6.700 ;
        RECT 15.950 5.950 16.950 6.550 ;
        RECT 13.450 5.700 16.550 6.300 ;
        RECT 3.700 5.950 14.050 6.550 ;
    END
  END b
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 2.350 13.550 3.050 16.250 ;
        RECT 0.000 13.750 18.750 16.250 ;
        RECT 5.750 13.550 6.450 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.200 7.200 13.200 7.800 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 7.500 8.400 14.900 9.000 ;
        RECT 4.100 10.950 18.300 11.550 ;
        RECT 14.650 6.800 15.250 7.900 ;
        RECT 14.650 7.300 18.300 7.900 ;
        RECT 4.100 4.600 18.300 5.200 ;
  END 
END exor2_4

MACRO exor2_3
  CLASS  CORE ;
  FOREIGN exor2_3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.750 9.700 2.750 10.300 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 10.500 0.000 11.100 2.650 ;
        RECT 0.000 0.000 15.000 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 12.300 9.700 14.300 10.300 ;
    END
  END b
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 1.550 13.100 2.150 16.250 ;
        RECT 0.000 13.750 15.000 16.250 ;
        RECT 3.700 13.100 4.300 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.850 9.700 7.850 10.300 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 5.400 5.950 9.400 6.550 ;
        RECT 9.950 6.650 10.550 7.650 ;
        RECT 0.450 7.050 10.550 7.650 ;
        RECT 5.400 3.150 12.950 3.750 ;
  END 
END exor2_3

MACRO exor2_2
  CLASS  CORE ;
  FOREIGN exor2_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.150 5.900 3.150 6.550 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 12.500 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.050 8.450 11.050 9.050 ;
    END
  END b
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 9.650 13.600 10.250 16.250 ;
        RECT 0.000 13.750 12.500 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.300 8.450 7.400 9.050 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 4.550 6.500 8.550 7.100 ;
  END 
END exor2_2

MACRO exor2_1
  CLASS  CORE ;
  FOREIGN exor2_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.450 7.200 7.450 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 10.000 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.750 8.450 9.750 9.050 ;
    END
  END b
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 10.000 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.400 8.450 6.150 10.300 ;
        RECT 3.450 9.700 6.150 10.300 ;
    END
  END x
END exor2_1

MACRO exnor3_5
  CLASS  CORE ;
  FOREIGN exnor3_5 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 21.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.950 7.200 2.950 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 2.150 0.000 2.750 2.800 ;
        RECT 0.000 0.000 21.250 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.950 5.950 3.950 6.550 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.300 5.950 10.300 6.550 ;
    END
  END c
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 2.100 13.500 2.800 16.250 ;
        RECT 0.000 13.750 21.250 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 17.400 8.450 18.100 10.150 ;
        RECT 17.400 8.450 19.150 9.150 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 0.450 4.700 5.050 5.300 ;
        RECT 4.450 4.700 5.050 7.800 ;
        RECT 4.350 7.200 5.550 7.800 ;
        RECT 4.350 7.200 4.950 9.050 ;
        RECT 0.450 8.450 4.950 9.050 ;
        RECT 8.550 8.450 9.150 10.150 ;
        RECT 3.850 9.550 9.150 10.150 ;
        RECT 5.550 5.950 6.700 6.550 ;
        RECT 6.100 7.200 11.250 7.800 ;
        RECT 6.100 5.950 6.700 9.050 ;
        RECT 5.550 8.450 6.700 9.050 ;
        RECT 15.350 8.500 15.950 10.150 ;
        RECT 10.650 9.550 15.950 10.150 ;
        RECT 12.350 5.950 13.500 6.550 ;
        RECT 12.900 7.150 19.350 7.850 ;
        RECT 12.900 5.950 13.500 9.050 ;
        RECT 12.350 8.450 13.500 9.050 ;
  END 
END exnor3_5

MACRO exnor3_4
  CLASS  CORE ;
  FOREIGN exnor3_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 20.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.850 7.200 2.850 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 2.150 0.000 2.750 2.800 ;
        RECT 0.000 0.000 20.000 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.850 5.950 3.850 6.550 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.400 5.950 10.400 6.550 ;
    END
  END c
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 2.100 13.500 2.800 16.250 ;
        RECT 0.000 13.750 20.000 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 17.200 8.450 19.200 9.050 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 0.450 4.700 4.950 5.300 ;
        RECT 4.350 7.200 5.550 7.800 ;
        RECT 4.350 4.700 4.950 9.050 ;
        RECT 0.450 8.450 4.950 9.050 ;
        RECT 8.550 8.450 9.150 10.150 ;
        RECT 3.850 9.550 9.150 10.150 ;
        RECT 5.550 6.100 6.700 6.700 ;
        RECT 6.100 7.200 11.250 7.800 ;
        RECT 6.100 6.100 6.700 9.050 ;
        RECT 5.550 8.450 6.700 9.050 ;
        RECT 15.350 8.500 15.950 10.150 ;
        RECT 10.650 9.550 15.950 10.150 ;
        RECT 12.350 7.150 19.150 7.850 ;
        RECT 12.350 5.950 12.950 9.050 ;
  END 
END exnor3_4

MACRO exnor3_3
  CLASS  CORE ;
  FOREIGN exnor3_3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 18.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.850 7.200 2.900 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 2.150 0.000 2.750 2.800 ;
        RECT 0.000 0.000 18.750 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.150 5.950 3.150 6.550 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.150 5.950 10.150 6.550 ;
    END
  END c
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 2.100 13.500 2.800 16.250 ;
        RECT 0.000 13.750 18.750 16.250 ;
        RECT 15.750 13.300 16.350 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 17.400 5.150 18.100 9.050 ;
        RECT 17.200 8.450 18.100 9.050 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 0.450 4.700 4.950 5.300 ;
        RECT 4.350 7.200 5.550 7.800 ;
        RECT 4.350 4.700 4.950 9.050 ;
        RECT 0.450 8.450 4.950 9.050 ;
        RECT 8.550 8.450 9.150 10.150 ;
        RECT 3.850 9.550 9.150 10.150 ;
        RECT 5.550 5.950 6.700 6.550 ;
        RECT 6.100 7.200 11.250 7.800 ;
        RECT 6.100 5.950 6.700 9.050 ;
        RECT 5.550 8.450 6.700 9.050 ;
        RECT 10.650 4.700 11.250 10.150 ;
        RECT 15.350 8.350 15.950 10.150 ;
        RECT 10.650 9.550 15.950 10.150 ;
        RECT 12.350 6.250 16.500 6.850 ;
        RECT 12.350 5.950 12.950 9.050 ;
  END 
END exnor3_3

MACRO exnor3_2
  CLASS  CORE ;
  FOREIGN exnor3_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 17.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.350 8.450 2.600 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 1.050 0.000 1.650 2.800 ;
        RECT 0.000 0.000 17.500 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.450 7.200 4.200 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.450 5.000 9.050 6.550 ;
        RECT 8.450 5.950 9.650 6.550 ;
    END
  END c
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.950 13.550 1.700 16.250 ;
        RECT 0.000 13.750 17.500 16.250 ;
        RECT 6.100 13.550 6.800 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 16.350 7.250 16.950 9.050 ;
        RECT 15.850 8.450 16.950 9.050 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 2.750 4.700 7.850 5.300 ;
        RECT 7.250 4.700 7.850 5.950 ;
        RECT 9.550 4.700 14.850 5.300 ;
        RECT 4.450 5.950 5.600 6.550 ;
        RECT 14.250 4.700 14.850 6.600 ;
        RECT 10.450 4.700 11.050 7.850 ;
        RECT 9.550 7.250 11.050 7.850 ;
        RECT 5.000 5.950 5.600 9.050 ;
        RECT 9.550 7.250 10.150 9.050 ;
        RECT 4.450 8.450 10.150 9.050 ;
        RECT 11.800 7.450 15.350 8.050 ;
        RECT 11.800 6.250 12.400 9.050 ;
        RECT 11.250 8.450 12.400 9.050 ;
  END 
END exnor3_2

MACRO exnor3_1
  CLASS  CORE ;
  FOREIGN exnor3_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 17.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.350 8.450 2.350 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 1.000 0.000 1.600 2.800 ;
        RECT 0.000 0.000 17.500 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.850 5.950 2.850 6.550 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.600 5.950 9.600 6.550 ;
    END
  END c
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.950 13.550 1.650 16.250 ;
        RECT 0.000 13.750 17.500 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 15.950 7.050 16.550 9.050 ;
        RECT 15.950 8.450 16.950 9.050 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 2.700 4.700 6.550 5.300 ;
        RECT 5.950 4.700 6.550 7.800 ;
        RECT 5.950 7.200 8.000 7.800 ;
        RECT 9.500 4.700 14.600 5.300 ;
        RECT 14.000 4.700 14.600 6.700 ;
        RECT 4.400 5.950 5.000 9.050 ;
        RECT 10.100 4.700 10.700 9.050 ;
        RECT 4.400 8.450 10.700 9.050 ;
        RECT 11.200 5.950 11.800 9.050 ;
        RECT 11.200 8.450 15.350 9.050 ;
  END 
END exnor3_1

MACRO exnor2_8
  CLASS  CORE ;
  FOREIGN exnor2_8 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 30.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.150 8.450 3.150 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 2.100 0.000 2.800 2.700 ;
        RECT 0.000 0.000 30.000 2.500 ;
        RECT 19.100 0.000 19.800 2.700 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.700 5.950 23.500 6.550 ;
    END
  END b
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 2.100 13.550 2.800 16.250 ;
        RECT 0.000 13.750 30.000 16.250 ;
        RECT 25.900 13.500 26.600 16.250 ;
        RECT 19.050 13.500 19.800 16.250 ;
        RECT 5.500 13.550 6.200 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.950 9.700 16.350 10.300 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 3.800 4.750 14.650 5.350 ;
        RECT 7.250 7.200 28.250 7.800 ;
        RECT 3.850 8.450 29.550 9.050 ;
  END 
END exnor2_8

MACRO exnor2_6
  CLASS  CORE ;
  FOREIGN exnor2_6 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 23.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.150 8.450 3.150 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 2.100 0.000 2.800 2.700 ;
        RECT 0.000 0.000 23.750 2.500 ;
        RECT 20.800 0.000 21.500 2.700 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.200 5.950 9.050 6.550 ;
        RECT 8.450 5.750 16.600 6.350 ;
    END
  END b
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 2.100 13.550 2.800 16.250 ;
        RECT 0.000 13.750 23.750 16.250 ;
        RECT 19.100 13.500 19.800 16.250 ;
        RECT 15.700 13.500 16.400 16.250 ;
        RECT 5.500 13.550 6.200 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.950 9.700 12.950 10.300 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 3.850 8.450 18.050 9.050 ;
        RECT 10.650 6.950 21.450 7.550 ;
        RECT 10.650 6.850 11.250 7.800 ;
        RECT 7.250 7.200 11.250 7.800 ;
  END 
END exnor2_6

MACRO exnor2_5
  CLASS  CORE ;
  FOREIGN exnor2_5 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 22.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.150 5.950 3.150 6.550 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 22.500 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.150 5.950 17.300 6.550 ;
    END
  END b
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 15.700 13.500 16.400 16.250 ;
        RECT 0.000 13.750 22.500 16.250 ;
        RECT 19.100 13.500 19.800 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.950 4.700 12.950 5.300 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 3.850 10.950 18.050 11.550 ;
        RECT 7.250 8.000 21.450 8.600 ;
  END 
END exnor2_5

MACRO exnor2_4
  CLASS  CORE ;
  FOREIGN exnor2_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 18.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.800 7.000 2.450 7.900 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 15.950 0.000 16.650 2.700 ;
        RECT 0.000 0.000 18.750 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.700 5.700 4.700 6.700 ;
        RECT 15.750 5.700 16.950 6.600 ;
        RECT 3.700 5.700 16.950 6.300 ;
    END
  END b
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 2.350 13.550 3.050 16.250 ;
        RECT 0.000 13.750 18.750 16.250 ;
        RECT 5.750 13.550 6.450 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.200 7.200 13.200 7.800 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 7.500 8.450 14.900 9.050 ;
        RECT 4.100 10.950 18.300 11.550 ;
        RECT 14.450 6.800 15.050 7.800 ;
        RECT 14.450 7.200 18.300 7.800 ;
        RECT 4.100 4.600 18.350 5.200 ;
  END 
END exnor2_4

MACRO exnor2_3
  CLASS  CORE ;
  FOREIGN exnor2_3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 10.000 6.650 10.600 7.800 ;
        RECT 0.750 7.200 10.600 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 10.500 0.000 11.100 2.650 ;
        RECT 0.000 0.000 15.000 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 12.400 9.700 14.400 10.300 ;
    END
  END b
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 1.550 13.100 2.150 16.250 ;
        RECT 0.000 13.750 15.000 16.250 ;
        RECT 3.700 13.100 4.300 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.900 9.700 7.900 10.300 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 5.400 5.950 9.400 6.550 ;
        RECT 5.400 3.150 12.950 3.750 ;
  END 
END exnor2_3

MACRO exnor2_2
  CLASS  CORE ;
  FOREIGN exnor2_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.150 5.950 3.150 6.550 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 12.500 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.700 8.450 11.700 9.050 ;
    END
  END b
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 9.650 13.600 10.250 16.250 ;
        RECT 0.000 13.750 12.500 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.400 8.450 7.400 9.050 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 4.550 6.500 8.600 7.100 ;
  END 
END exnor2_2

MACRO exnor2_1
  CLASS  CORE ;
  FOREIGN exnor2_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.650 7.200 7.900 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 10.000 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.600 4.700 9.600 5.300 ;
    END
  END b
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 10.000 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.150 5.950 6.450 6.550 ;
    END
  END x
END exnor2_1

MACRO dffpt_8
  CLASS  CORE ;
  FOREIGN dffpt_8 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 30.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 24.350 8.450 26.350 9.050 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 2.250 0.000 2.850 2.800 ;
        RECT 0.000 0.000 30.000 2.500 ;
        RECT 9.300 0.000 9.900 2.800 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.550 7.200 4.550 7.800 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 1.000 13.500 1.600 16.250 ;
        RECT 0.000 13.750 30.000 16.250 ;
        RECT 20.100 13.450 20.700 16.250 ;
    END
  END vdd!
  PIN setb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.400 5.950 2.400 6.550 ;
    END
  END setb
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 20.400 8.450 22.900 9.050 ;
    END
  END qb
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 27.300 4.700 29.350 5.300 ;
    END
  END ck
  OBS 
      LAYER Metal1 ;
        RECT 5.050 4.700 6.250 5.300 ;
        RECT 5.050 4.700 5.650 10.150 ;
        RECT 5.050 9.550 6.750 10.150 ;
        RECT 6.150 5.950 15.000 6.550 ;
        RECT 6.150 5.950 6.750 9.050 ;
        RECT 6.150 8.450 12.300 9.050 ;
        RECT 10.400 9.600 11.000 10.300 ;
        RECT 10.400 9.700 19.000 10.300 ;
        RECT 12.500 4.700 24.500 5.300 ;
        RECT 14.750 7.050 15.350 7.800 ;
        RECT 7.250 7.200 29.200 7.800 ;
        RECT 7.250 7.200 7.850 7.950 ;
  END 
END dffpt_8

MACRO dffpt_6
  CLASS  CORE ;
  FOREIGN dffpt_6 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 28.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 22.750 9.700 25.350 10.300 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 2.250 0.000 2.850 2.800 ;
        RECT 0.000 0.000 28.750 2.500 ;
        RECT 22.550 0.000 23.150 2.650 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.100 7.200 4.100 7.800 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 22.550 13.450 23.150 16.250 ;
        RECT 0.000 13.750 28.750 16.250 ;
    END
  END vdd!
  PIN setb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.400 5.950 2.400 6.550 ;
    END
  END setb
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 17.850 8.450 19.850 9.050 ;
    END
  END qb
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 26.250 5.950 28.250 6.550 ;
    END
  END ck
  OBS 
      LAYER Metal1 ;
        RECT 4.600 4.700 6.350 5.300 ;
        RECT 4.600 4.700 5.200 10.300 ;
        RECT 4.600 9.700 6.350 10.300 ;
        RECT 5.700 5.950 14.800 6.550 ;
        RECT 5.700 5.950 6.300 8.950 ;
        RECT 5.700 8.350 11.600 8.950 ;
        RECT 9.700 9.500 10.300 10.250 ;
        RECT 9.700 9.650 21.450 10.250 ;
        RECT 16.500 7.100 22.750 7.700 ;
        RECT 16.500 7.100 17.100 8.950 ;
        RECT 12.350 8.350 17.100 8.950 ;
        RECT 15.400 6.000 24.500 6.600 ;
        RECT 23.900 6.000 24.500 7.800 ;
        RECT 15.400 6.000 16.000 7.800 ;
        RECT 6.800 7.200 16.000 7.800 ;
        RECT 23.900 7.200 28.300 7.800 ;
        RECT 6.800 7.200 7.400 7.850 ;
        RECT 14.200 7.200 14.800 7.850 ;
  END 
END dffpt_6

MACRO dffpt_4
  CLASS  CORE ;
  FOREIGN dffpt_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 27.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 22.850 7.200 24.850 7.800 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 27.500 2.500 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.850 8.450 4.850 9.050 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 27.500 16.250 ;
    END
  END vdd!
  PIN setb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 7.200 2.300 7.800 ;
    END
  END setb
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 19.250 5.950 21.250 6.550 ;
    END
  END qb
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.950 5.950 11.950 6.550 ;
    END
  END ck
  OBS 
      LAYER Metal1 ;
        RECT 6.200 6.050 7.500 6.650 ;
        RECT 6.200 6.050 6.800 7.950 ;
        RECT 5.350 7.350 6.800 7.950 ;
        RECT 5.350 7.350 5.950 10.150 ;
        RECT 5.350 9.550 7.550 10.150 ;
        RECT 12.650 6.250 18.200 6.850 ;
        RECT 7.600 7.150 8.200 7.950 ;
        RECT 12.650 6.250 13.250 7.950 ;
        RECT 7.600 7.350 13.300 7.950 ;
        RECT 17.600 6.250 18.200 7.950 ;
        RECT 14.350 7.350 14.950 9.050 ;
        RECT 6.650 8.450 19.250 9.050 ;
  END 
END dffpt_4

MACRO dffpt_3
  CLASS  CORE ;
  FOREIGN dffpt_3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 25.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 20.900 5.950 22.900 6.550 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 9.650 0.000 10.250 2.800 ;
        RECT 0.000 0.000 25.000 2.500 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.650 8.450 4.650 9.050 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 25.000 16.250 ;
    END
  END vdd!
  PIN setb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.550 7.200 2.550 7.800 ;
    END
  END setb
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 18.250 5.950 20.250 6.550 ;
    END
  END qb
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.650 5.950 11.650 6.550 ;
    END
  END ck
  OBS 
      LAYER Metal1 ;
        RECT 6.300 6.150 7.500 6.750 ;
        RECT 6.300 6.150 6.900 7.850 ;
        RECT 5.500 7.250 6.900 7.850 ;
        RECT 5.500 7.250 6.100 10.250 ;
        RECT 5.500 9.650 7.600 10.250 ;
        RECT 6.800 8.450 17.650 9.050 ;
        RECT 6.800 8.450 7.400 9.150 ;
        RECT 7.550 7.250 8.150 7.950 ;
        RECT 7.550 7.350 18.250 7.950 ;
  END 
END dffpt_3

MACRO dffpt_2
  CLASS  CORE ;
  FOREIGN dffpt_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 21.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 15.900 8.400 17.850 9.050 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 9.050 0.000 9.650 2.700 ;
        RECT 0.000 0.000 21.250 2.500 ;
        RECT 15.050 0.000 15.650 2.800 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.650 8.450 3.650 9.050 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 1.850 13.550 2.450 16.250 ;
        RECT 0.000 13.750 21.250 16.250 ;
        RECT 9.150 13.550 9.750 16.250 ;
    END
  END vdd!
  PIN setb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.850 5.950 2.850 6.550 ;
    END
  END setb
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 13.200 8.450 15.200 9.050 ;
    END
  END qb
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 18.500 8.450 20.500 9.050 ;
    END
  END ck
  OBS 
      LAYER Metal1 ;
        RECT 5.350 5.800 5.950 6.550 ;
        RECT 4.350 5.950 5.950 6.550 ;
        RECT 4.350 5.950 4.950 9.200 ;
        RECT 4.350 8.600 6.550 9.200 ;
        RECT 6.450 6.250 11.350 6.850 ;
        RECT 6.450 6.250 7.050 7.650 ;
        RECT 5.450 7.050 7.050 7.650 ;
        RECT 5.450 7.050 6.050 8.100 ;
        RECT 12.050 7.250 20.850 7.850 ;
        RECT 7.550 7.350 12.650 7.950 ;
  END 
END dffpt_2

MACRO dffpt_1
  CLASS  CORE ;
  FOREIGN dffpt_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 20.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 17.650 5.950 19.650 6.550 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 2.050 0.000 2.650 2.700 ;
        RECT 0.000 0.000 20.000 2.500 ;
        RECT 17.300 0.000 17.900 2.700 ;
        RECT 11.200 0.000 11.800 2.700 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.150 8.450 3.150 9.050 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 1.850 13.550 2.450 16.250 ;
        RECT 0.000 13.750 20.000 16.250 ;
        RECT 17.250 13.550 17.850 16.250 ;
        RECT 9.450 13.550 10.050 16.250 ;
    END
  END vdd!
  PIN setb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.800 5.950 2.800 6.550 ;
    END
  END setb
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 17.200 8.450 19.200 9.050 ;
    END
  END qb
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.550 3.450 10.550 4.050 ;
    END
  END ck
  OBS 
      LAYER Metal1 ;
        RECT 5.500 5.800 6.100 6.550 ;
        RECT 3.750 5.950 6.100 6.550 ;
        RECT 3.750 5.950 4.350 9.200 ;
        RECT 3.750 8.600 6.550 9.200 ;
        RECT 6.750 6.250 12.800 6.850 ;
        RECT 6.750 6.250 7.350 7.650 ;
        RECT 4.850 7.050 7.350 7.650 ;
        RECT 4.850 7.050 5.450 8.100 ;
        RECT 12.200 8.450 15.400 9.050 ;
        RECT 10.900 7.350 16.100 7.950 ;
        RECT 10.900 7.350 11.500 8.950 ;
        RECT 7.450 8.350 11.500 8.950 ;
  END 
END dffpt_1

MACRO dffps_8
  CLASS  CORE ;
  FOREIGN dffps_8 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 30.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN sb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.350 8.450 2.400 9.050 ;
    END
  END sb
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 18.250 8.450 22.750 9.050 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 19.950 0.000 20.550 2.800 ;
        RECT 0.000 0.000 30.000 2.500 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.100 5.950 3.100 6.550 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 19.950 13.450 20.550 16.250 ;
        RECT 0.000 13.750 30.000 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 24.200 9.700 26.200 10.300 ;
    END
  END qb
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 27.150 4.700 29.150 5.300 ;
    END
  END ck
  OBS 
      LAYER Metal1 ;
        RECT 3.650 4.700 5.200 5.300 ;
        RECT 3.650 4.700 4.250 10.300 ;
        RECT 3.650 9.700 4.900 10.300 ;
        RECT 4.750 6.250 13.700 6.850 ;
        RECT 4.750 6.250 5.350 9.050 ;
        RECT 4.750 8.450 10.500 9.050 ;
        RECT 8.600 9.550 9.200 10.250 ;
        RECT 8.600 9.650 17.550 10.250 ;
        RECT 11.200 4.700 20.100 5.300 ;
        RECT 23.750 5.700 24.350 6.550 ;
        RECT 18.200 5.950 24.350 6.550 ;
        RECT 15.300 7.200 29.050 7.800 ;
        RECT 5.850 7.350 15.900 7.950 ;
        RECT 12.900 7.350 13.500 8.300 ;
  END 
END dffps_8

MACRO dffps_6
  CLASS  CORE ;
  FOREIGN dffps_6 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 27.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN sb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.300 8.450 2.300 9.050 ;
    END
  END sb
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 21.850 9.700 23.850 10.300 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 18.050 0.000 18.650 2.800 ;
        RECT 0.000 0.000 27.500 2.500 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.250 4.700 3.250 5.300 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 21.050 13.450 21.650 16.250 ;
        RECT 0.000 13.750 27.500 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 15.550 5.950 17.550 6.550 ;
    END
  END qb
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 24.950 5.950 26.950 6.550 ;
    END
  END ck
  OBS 
      LAYER Metal1 ;
        RECT 2.550 6.000 3.400 6.600 ;
        RECT 2.800 6.000 3.400 10.300 ;
        RECT 2.450 9.650 3.400 10.300 ;
        RECT 3.900 4.700 4.950 5.300 ;
        RECT 3.900 4.700 4.500 10.150 ;
        RECT 3.900 9.550 5.600 10.150 ;
        RECT 12.800 6.050 13.400 6.750 ;
        RECT 5.050 6.150 13.400 6.750 ;
        RECT 5.050 6.150 5.650 9.050 ;
        RECT 7.250 8.350 10.050 8.950 ;
        RECT 5.000 8.450 7.850 9.050 ;
        RECT 6.300 4.950 14.900 5.550 ;
        RECT 6.300 4.950 6.900 5.650 ;
        RECT 14.300 4.950 14.900 6.650 ;
        RECT 8.450 9.500 9.050 10.250 ;
        RECT 8.450 9.650 19.950 10.250 ;
        RECT 18.850 5.950 21.650 6.550 ;
        RECT 10.850 8.450 24.650 9.050 ;
        RECT 6.150 7.250 26.900 7.850 ;
        RECT 6.150 7.250 6.750 7.950 ;
        RECT 12.800 7.250 13.400 7.950 ;
  END 
END dffps_6

MACRO dffps_4
  CLASS  CORE ;
  FOREIGN dffps_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 22.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN sb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 7.200 2.250 7.800 ;
    END
  END sb
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 16.050 9.700 18.050 10.300 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 11.000 0.000 11.600 2.650 ;
        RECT 0.000 0.000 22.500 2.500 ;
        RECT 15.600 0.000 16.200 3.750 ;
        RECT 13.200 0.000 13.800 2.650 ;
        RECT 12.100 0.000 12.700 2.650 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.650 9.700 2.950 10.300 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 22.500 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 13.350 9.700 15.350 10.300 ;
    END
  END qb
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 20.250 5.950 22.250 6.550 ;
    END
  END ck
  OBS 
      LAYER Metal1 ;
        RECT 4.000 5.850 4.600 7.750 ;
        RECT 3.450 7.150 4.050 10.300 ;
        RECT 3.450 9.700 5.650 10.300 ;
        RECT 5.550 7.150 10.450 7.750 ;
        RECT 9.850 7.150 10.450 8.100 ;
        RECT 10.050 5.850 11.550 6.450 ;
        RECT 10.950 7.350 16.350 7.950 ;
        RECT 10.950 5.850 11.550 9.250 ;
        RECT 12.050 5.850 19.750 6.450 ;
        RECT 19.150 5.850 19.750 7.050 ;
        RECT 4.550 8.250 9.350 8.850 ;
        RECT 20.450 8.000 21.050 9.050 ;
        RECT 12.250 8.450 21.050 9.050 ;
        RECT 8.750 8.250 9.350 10.400 ;
        RECT 12.250 8.450 12.850 10.400 ;
        RECT 8.750 9.800 12.850 10.400 ;
  END 
END dffps_4

MACRO dffps_3
  CLASS  CORE ;
  FOREIGN dffps_3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 22.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN sb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 7.200 2.250 7.800 ;
    END
  END sb
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 16.800 10.950 18.800 11.550 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 22.500 2.500 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.150 9.600 1.750 11.550 ;
        RECT 1.150 10.850 2.900 11.550 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 22.500 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 13.300 10.950 15.300 11.550 ;
    END
  END qb
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 21.650 6.950 22.250 10.300 ;
        RECT 20.750 9.600 22.250 10.300 ;
    END
  END ck
  OBS 
      LAYER Metal1 ;
        RECT 3.100 6.050 4.600 6.650 ;
        RECT 3.100 6.050 3.700 10.100 ;
        RECT 3.100 9.500 5.600 10.100 ;
        RECT 5.600 7.150 10.600 7.750 ;
        RECT 9.650 5.850 11.700 6.450 ;
        RECT 15.850 7.350 16.450 8.900 ;
        RECT 11.100 8.300 16.450 8.900 ;
        RECT 11.100 5.850 11.700 9.250 ;
        RECT 12.200 5.850 19.750 6.450 ;
        RECT 12.200 5.850 12.800 7.750 ;
        RECT 19.150 5.850 19.750 7.950 ;
        RECT 20.350 5.850 21.150 6.450 ;
        RECT 4.400 8.250 9.500 8.850 ;
        RECT 20.350 5.850 20.950 9.100 ;
        RECT 19.250 8.500 20.950 9.100 ;
        RECT 8.900 8.250 9.500 10.350 ;
        RECT 12.500 9.400 19.850 10.000 ;
        RECT 19.250 8.500 19.850 10.000 ;
        RECT 8.900 9.750 13.100 10.350 ;
  END 
END dffps_3

MACRO dffps_2
  CLASS  CORE ;
  FOREIGN dffps_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 21.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN sb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 8.450 2.250 9.050 ;
    END
  END sb
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 15.450 5.950 17.450 6.550 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 1.000 0.000 1.600 2.700 ;
        RECT 0.000 0.000 21.250 2.500 ;
        RECT 14.500 0.000 15.100 3.800 ;
        RECT 6.100 0.000 6.700 2.800 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.000 5.950 3.000 6.550 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 1.000 13.550 1.600 16.250 ;
        RECT 0.000 13.750 21.250 16.250 ;
        RECT 14.500 13.550 15.100 16.250 ;
        RECT 6.200 13.550 6.800 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 12.600 5.950 14.600 6.550 ;
    END
  END qb
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 18.950 7.200 20.950 7.800 ;
    END
  END ck
  OBS 
      LAYER Metal1 ;
        RECT 5.700 8.500 9.550 9.100 ;
        RECT 8.950 8.500 9.550 9.200 ;
        RECT 4.100 5.200 9.750 5.800 ;
        RECT 4.100 5.200 4.700 6.600 ;
        RECT 3.500 6.000 4.100 9.200 ;
        RECT 3.500 8.600 5.200 9.200 ;
        RECT 5.700 6.300 12.100 6.900 ;
        RECT 11.500 5.200 12.100 7.950 ;
        RECT 11.500 7.350 18.450 7.950 ;
        RECT 4.600 7.400 10.650 8.000 ;
        RECT 4.600 7.400 5.200 8.100 ;
        RECT 10.050 7.400 10.650 9.050 ;
        RECT 10.050 8.450 19.800 9.050 ;
  END 
END dffps_2

MACRO dffps_1
  CLASS  CORE ;
  FOREIGN dffps_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 21.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN sb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.950 7.500 1.550 9.050 ;
        RECT 0.250 8.450 1.550 9.050 ;
    END
  END sb
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 15.250 5.950 17.250 6.550 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 1.000 0.000 1.600 2.700 ;
        RECT 0.000 0.000 21.250 2.500 ;
        RECT 17.300 0.000 17.900 2.600 ;
        RECT 14.300 0.000 14.900 3.750 ;
        RECT 6.100 0.000 6.700 2.800 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.000 4.700 1.700 6.550 ;
        RECT 1.000 4.700 2.900 5.400 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 1.000 13.550 1.600 16.250 ;
        RECT 0.000 13.750 21.250 16.250 ;
        RECT 6.350 13.550 6.950 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 12.600 5.950 14.600 6.550 ;
    END
  END qb
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 18.950 7.200 20.950 7.800 ;
    END
  END ck
  OBS 
      LAYER Metal1 ;
        RECT 5.700 8.500 9.550 9.100 ;
        RECT 8.950 8.500 9.550 9.200 ;
        RECT 4.100 5.200 9.750 5.800 ;
        RECT 4.100 5.200 4.700 6.600 ;
        RECT 2.350 6.000 4.700 6.600 ;
        RECT 2.350 6.000 2.950 9.200 ;
        RECT 2.350 8.600 5.200 9.200 ;
        RECT 5.700 6.300 12.100 6.900 ;
        RECT 11.500 5.200 12.100 7.950 ;
        RECT 11.500 7.350 18.450 7.950 ;
        RECT 4.600 7.400 10.650 8.000 ;
        RECT 3.500 7.500 5.200 8.100 ;
        RECT 10.050 7.400 10.650 9.050 ;
        RECT 10.050 8.450 19.800 9.050 ;
  END 
END dffps_1

MACRO dffprs_8
  CLASS  CORE ;
  FOREIGN dffprs_8 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 31.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN sb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 10.550 9.600 11.150 10.450 ;
        RECT 10.550 9.850 19.050 10.450 ;
        RECT 18.450 8.450 19.050 10.450 ;
    END
  END sb
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 24.250 9.700 26.350 10.300 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.500 0.000 1.100 2.800 ;
        RECT 0.000 0.000 31.250 2.500 ;
        RECT 20.100 0.000 20.700 2.800 ;
        RECT 11.400 0.000 12.000 2.800 ;
        RECT 9.700 0.000 10.300 2.800 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.950 7.500 1.550 9.050 ;
        RECT 0.300 8.450 1.550 9.050 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 10.200 13.450 10.800 16.250 ;
        RECT 0.000 13.750 31.250 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 21.200 9.700 23.350 10.300 ;
    END
  END qb
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 28.900 7.200 30.900 7.800 ;
    END
  END ck
  PIN rb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.200 5.950 2.800 10.300 ;
        RECT 8.950 5.950 9.550 6.900 ;
        RECT 0.350 5.950 9.550 6.550 ;
        RECT 2.200 9.700 6.300 10.300 ;
    END
  END rb
  OBS 
      LAYER Metal1 ;
        RECT 11.650 7.350 14.200 7.950 ;
        RECT 5.500 4.700 24.500 5.300 ;
        RECT 17.050 7.250 28.300 7.850 ;
        RECT 4.600 8.500 13.150 9.100 ;
        RECT 17.050 7.250 17.650 9.350 ;
        RECT 12.550 8.750 17.650 9.350 ;
        RECT 8.300 8.500 8.900 9.800 ;
        RECT 10.150 6.000 29.600 6.600 ;
        RECT 10.150 6.000 10.750 8.000 ;
        RECT 3.500 7.400 10.750 8.000 ;
        RECT 15.450 6.000 16.050 8.250 ;
  END 
END dffprs_8

MACRO dffprs_6
  CLASS  CORE ;
  FOREIGN dffprs_6 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 30.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN sb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 18.450 8.450 19.050 10.300 ;
        RECT 10.850 9.700 19.050 10.300 ;
    END
  END sb
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 23.800 9.700 25.800 10.300 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.500 0.000 1.100 2.800 ;
        RECT 0.000 0.000 30.000 2.500 ;
        RECT 19.550 0.000 20.150 2.800 ;
        RECT 12.400 0.000 13.000 2.800 ;
        RECT 10.450 0.000 11.050 2.800 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.950 7.500 1.550 9.050 ;
        RECT 0.300 8.450 1.550 9.050 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 9.300 13.450 9.900 16.250 ;
        RECT 0.000 13.750 30.000 16.250 ;
        RECT 13.850 13.450 14.450 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 20.650 9.700 22.650 10.300 ;
    END
  END qb
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 27.650 7.200 29.650 7.800 ;
    END
  END ck
  PIN rb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.200 5.950 2.800 10.300 ;
        RECT 9.600 5.950 10.200 6.900 ;
        RECT 9.150 5.950 10.200 6.650 ;
        RECT 0.350 5.950 10.200 6.550 ;
        RECT 2.200 9.700 5.800 10.300 ;
    END
  END rb
  OBS 
      LAYER Metal1 ;
        RECT 12.150 7.350 14.450 7.950 ;
        RECT 5.550 4.700 23.950 5.300 ;
        RECT 16.800 7.250 27.100 7.850 ;
        RECT 16.800 7.250 17.400 9.100 ;
        RECT 4.800 8.500 17.400 9.100 ;
        RECT 10.800 6.000 28.350 6.600 ;
        RECT 15.700 6.000 16.300 7.850 ;
        RECT 10.800 6.000 11.400 8.000 ;
        RECT 3.500 7.400 11.400 8.000 ;
  END 
END dffprs_6

MACRO dffprs_4
  CLASS  CORE ;
  FOREIGN dffprs_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 27.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN sb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 14.100 9.550 14.700 10.300 ;
        RECT 14.100 9.700 16.050 10.300 ;
    END
  END sb
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 21.050 9.700 23.050 10.300 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 10.100 0.000 10.800 2.800 ;
        RECT 0.000 0.000 27.500 2.500 ;
        RECT 12.150 0.000 12.750 2.700 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.300 8.450 2.300 9.050 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 27.500 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 17.550 9.700 19.550 10.300 ;
    END
  END qb
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 26.650 6.700 27.250 10.300 ;
        RECT 25.950 9.700 27.250 10.300 ;
    END
  END ck
  PIN rb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.350 5.950 10.600 6.550 ;
        RECT 10.000 5.950 10.600 6.800 ;
    END
  END rb
  OBS 
      LAYER Metal1 ;
        RECT 10.250 9.800 13.400 10.400 ;
        RECT 5.950 4.600 16.450 5.200 ;
        RECT 21.000 6.750 21.600 7.400 ;
        RECT 15.700 6.800 21.600 7.400 ;
        RECT 19.600 5.600 24.700 6.200 ;
        RECT 11.600 5.700 20.250 6.300 ;
        RECT 24.100 5.600 24.700 7.050 ;
        RECT 4.650 7.150 5.250 7.950 ;
        RECT 11.600 5.700 12.200 7.950 ;
        RECT 4.650 7.350 12.200 7.950 ;
        RECT 7.900 7.350 8.500 8.850 ;
        RECT 25.400 5.450 26.300 6.100 ;
        RECT 17.300 7.900 17.900 9.050 ;
        RECT 25.400 5.450 26.000 9.050 ;
        RECT 9.000 8.450 26.000 9.050 ;
        RECT 9.000 8.450 9.600 9.950 ;
        RECT 3.250 9.350 9.600 9.950 ;
  END 
END dffprs_4

MACRO dffprs_3
  CLASS  CORE ;
  FOREIGN dffprs_3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 26.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN sb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 14.100 9.550 14.700 10.300 ;
        RECT 14.100 9.700 15.950 10.300 ;
    END
  END sb
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 20.550 9.700 22.550 10.300 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 10.450 0.000 11.050 2.800 ;
        RECT 0.000 0.000 26.250 2.500 ;
        RECT 12.150 0.000 12.750 2.700 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.300 8.450 2.300 9.050 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 15.950 13.550 16.550 16.250 ;
        RECT 0.000 13.750 26.250 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 17.050 9.700 19.050 10.300 ;
    END
  END qb
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 24.700 4.700 26.000 5.300 ;
        RECT 25.400 4.700 26.000 8.200 ;
    END
  END ck
  PIN rb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.350 5.950 10.200 6.550 ;
        RECT 9.150 5.950 10.200 6.800 ;
    END
  END rb
  OBS 
      LAYER Metal1 ;
        RECT 10.300 9.550 13.400 10.150 ;
        RECT 6.250 4.600 16.050 5.200 ;
        RECT 15.450 8.450 20.350 9.050 ;
        RECT 11.600 5.700 23.200 6.300 ;
        RECT 22.600 5.700 23.200 7.250 ;
        RECT 4.650 7.150 8.500 7.800 ;
        RECT 11.600 5.700 12.200 7.900 ;
        RECT 7.900 7.300 12.200 7.900 ;
        RECT 7.900 7.150 8.500 8.700 ;
        RECT 14.050 6.950 21.650 7.550 ;
        RECT 21.050 6.950 21.650 8.400 ;
        RECT 21.050 7.800 24.900 8.400 ;
        RECT 24.300 6.250 24.900 9.400 ;
        RECT 14.050 6.950 14.650 9.050 ;
        RECT 9.200 8.450 14.650 9.050 ;
        RECT 24.300 8.800 25.050 9.400 ;
        RECT 3.900 9.350 9.800 9.950 ;
        RECT 9.200 8.450 9.800 9.950 ;
        RECT 3.250 9.550 4.500 10.150 ;
  END 
END dffprs_3

MACRO dffprs_2
  CLASS  CORE ;
  FOREIGN dffprs_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 26.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN sb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 13.450 9.700 15.450 10.300 ;
    END
  END sb
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 20.250 9.700 22.250 10.300 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 10.100 0.000 10.700 2.700 ;
        RECT 0.000 0.000 26.250 2.500 ;
        RECT 12.550 0.000 13.150 2.700 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.600 8.450 2.600 9.050 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 10.600 13.550 11.200 16.250 ;
        RECT 0.000 13.750 26.250 16.250 ;
        RECT 14.050 13.550 14.650 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 16.850 9.700 18.850 10.300 ;
    END
  END qb
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 25.300 6.400 25.900 7.800 ;
        RECT 24.500 7.200 25.900 7.800 ;
    END
  END ck
  PIN rb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.350 5.950 5.400 6.550 ;
    END
  END rb
  OBS 
      LAYER Metal1 ;
        RECT 5.400 3.450 11.850 4.050 ;
        RECT 10.100 9.750 12.950 10.350 ;
        RECT 11.250 7.350 20.050 7.950 ;
        RECT 7.650 7.550 11.850 8.150 ;
        RECT 7.650 7.550 8.250 8.850 ;
        RECT 5.900 8.250 8.250 8.850 ;
        RECT 10.150 6.250 23.100 6.850 ;
        RECT 5.900 6.450 10.750 7.050 ;
        RECT 5.900 6.450 6.500 7.750 ;
        RECT 3.500 7.150 6.500 7.750 ;
        RECT 22.500 6.250 23.100 7.800 ;
        RECT 12.350 8.450 24.950 9.050 ;
        RECT 9.000 8.650 12.950 9.250 ;
        RECT 9.000 8.650 9.600 9.950 ;
        RECT 3.500 9.350 9.600 9.950 ;
  END 
END dffprs_2

MACRO dffprs_1
  CLASS  CORE ;
  FOREIGN dffprs_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 26.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN sb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 13.450 9.700 15.450 10.300 ;
    END
  END sb
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 20.250 9.700 22.250 10.300 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 10.100 0.000 10.700 2.700 ;
        RECT 0.000 0.000 26.250 2.500 ;
        RECT 12.550 0.000 13.150 2.700 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.600 8.450 2.600 9.050 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 10.600 13.550 11.200 16.250 ;
        RECT 0.000 13.750 26.250 16.250 ;
        RECT 14.050 13.550 14.650 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 16.850 9.700 18.850 10.300 ;
    END
  END qb
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 24.000 7.200 26.000 7.800 ;
    END
  END ck
  PIN rb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.350 5.950 5.400 6.550 ;
    END
  END rb
  OBS 
      LAYER Metal1 ;
        RECT 5.400 3.450 11.850 4.050 ;
        RECT 10.100 9.750 12.950 10.350 ;
        RECT 11.250 7.350 20.250 7.950 ;
        RECT 7.650 7.550 11.850 8.150 ;
        RECT 7.650 7.550 8.250 8.850 ;
        RECT 5.900 8.250 8.250 8.850 ;
        RECT 10.150 6.250 23.300 6.850 ;
        RECT 5.900 6.450 10.750 7.050 ;
        RECT 5.900 6.450 6.500 7.750 ;
        RECT 3.500 7.150 6.500 7.750 ;
        RECT 22.700 6.250 23.300 7.800 ;
        RECT 12.350 8.450 24.600 9.050 ;
        RECT 9.000 8.650 12.950 9.250 ;
        RECT 9.000 8.650 9.600 9.950 ;
        RECT 3.500 9.350 9.600 9.950 ;
  END 
END dffprs_1

MACRO dffpr_8
  CLASS  CORE ;
  FOREIGN dffpr_8 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 30.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 18.450 9.700 22.450 10.300 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 17.150 0.000 17.750 2.800 ;
        RECT 0.000 0.000 30.000 2.500 ;
        RECT 20.150 0.000 20.750 2.800 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.100 5.950 3.100 6.550 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 7.950 13.450 8.550 16.250 ;
        RECT 0.000 13.750 30.000 16.250 ;
        RECT 26.950 13.450 27.550 16.250 ;
        RECT 20.150 13.450 20.750 16.250 ;
        RECT 15.450 13.450 16.050 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 24.400 8.450 26.400 9.050 ;
    END
  END qb
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 27.350 4.700 29.450 5.300 ;
    END
  END ck
  PIN rb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.300 8.450 2.300 9.050 ;
    END
  END rb
  OBS 
      LAYER Metal1 ;
        RECT 4.000 6.250 5.000 6.850 ;
        RECT 4.000 6.250 4.600 10.150 ;
        RECT 4.000 9.550 5.850 10.150 ;
        RECT 12.750 6.050 13.350 6.850 ;
        RECT 5.500 6.250 13.350 6.850 ;
        RECT 5.500 6.250 6.100 9.050 ;
        RECT 5.400 8.450 10.950 9.050 ;
        RECT 8.250 4.950 15.450 5.550 ;
        RECT 8.250 4.950 8.850 5.750 ;
        RECT 14.850 4.950 15.450 6.850 ;
        RECT 9.050 9.550 9.650 10.250 ;
        RECT 9.050 9.650 17.750 10.250 ;
        RECT 11.650 8.450 21.150 9.050 ;
        RECT 18.850 5.300 24.550 5.900 ;
        RECT 16.500 7.200 29.250 7.800 ;
        RECT 6.800 7.350 17.100 7.950 ;
  END 
END dffpr_8

MACRO dffpr_6
  CLASS  CORE ;
  FOREIGN dffpr_6 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 27.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 22.100 9.700 24.100 10.300 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 16.600 0.000 17.200 2.800 ;
        RECT 0.000 0.000 27.500 2.500 ;
        RECT 24.700 0.000 25.300 2.800 ;
        RECT 21.300 0.000 21.900 2.800 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.950 5.950 2.950 6.550 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 7.400 13.450 8.000 16.250 ;
        RECT 0.000 13.750 27.500 16.250 ;
        RECT 21.300 13.450 21.900 16.250 ;
        RECT 18.300 13.450 18.900 16.250 ;
        RECT 14.900 13.450 15.500 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 16.850 5.950 18.900 6.550 ;
    END
  END qb
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 25.000 4.700 27.000 5.300 ;
    END
  END ck
  PIN rb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.350 8.450 2.350 9.050 ;
    END
  END rb
  OBS 
      LAYER Metal1 ;
        RECT 3.550 6.250 4.850 6.850 ;
        RECT 3.550 6.250 4.150 10.150 ;
        RECT 3.550 9.550 5.350 10.150 ;
        RECT 5.350 6.250 13.200 6.850 ;
        RECT 5.350 6.250 5.950 9.050 ;
        RECT 4.650 8.450 10.800 9.050 ;
        RECT 7.850 5.150 15.100 5.750 ;
        RECT 14.500 5.150 15.100 6.600 ;
        RECT 8.500 9.550 9.100 10.250 ;
        RECT 8.500 9.650 20.200 10.250 ;
        RECT 11.300 8.450 24.900 9.050 ;
        RECT 6.450 7.350 27.100 7.950 ;
  END 
END dffpr_6

MACRO dffpr_4
  CLASS  CORE ;
  FOREIGN dffpr_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 22.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 16.050 5.950 18.050 6.550 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 22.500 2.500 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.800 5.950 2.900 6.550 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 22.500 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 12.550 9.700 14.550 10.300 ;
    END
  END qb
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 21.550 6.850 22.150 10.300 ;
        RECT 20.750 9.700 22.150 10.300 ;
    END
  END ck
  PIN rb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 8.450 2.250 9.050 ;
    END
  END rb
  OBS 
      LAYER Metal1 ;
        RECT 4.000 6.100 10.500 6.700 ;
        RECT 4.000 6.100 4.600 7.800 ;
        RECT 3.000 7.200 4.600 7.800 ;
        RECT 3.000 7.200 3.600 10.300 ;
        RECT 3.000 9.700 5.850 10.300 ;
        RECT 12.600 6.200 13.200 7.950 ;
        RECT 19.300 6.450 19.900 7.950 ;
        RECT 5.600 7.350 19.900 7.950 ;
        RECT 5.600 7.350 6.200 8.100 ;
        RECT 20.400 4.700 21.300 5.300 ;
        RECT 4.100 8.300 4.700 9.200 ;
        RECT 7.500 8.450 21.000 9.050 ;
        RECT 20.400 4.700 21.000 9.050 ;
        RECT 4.100 8.600 8.100 9.200 ;
  END 
END dffpr_4

MACRO dffpr_3
  CLASS  CORE ;
  FOREIGN dffpr_3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 22.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 16.300 5.950 18.300 6.550 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 22.500 2.500 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.100 5.950 3.400 6.550 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 22.500 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 13.300 9.700 15.300 10.300 ;
    END
  END qb
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 21.550 5.250 22.150 6.550 ;
        RECT 20.850 5.950 22.150 6.550 ;
    END
  END ck
  PIN rb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 8.450 2.250 9.050 ;
    END
  END rb
  OBS 
      LAYER Metal1 ;
        RECT 4.400 6.100 10.350 6.700 ;
        RECT 4.400 6.100 5.000 7.700 ;
        RECT 3.500 7.100 5.000 7.700 ;
        RECT 3.500 7.100 4.100 10.300 ;
        RECT 3.500 9.700 5.100 10.300 ;
        RECT 12.550 6.350 13.150 7.950 ;
        RECT 6.000 7.350 19.750 7.950 ;
        RECT 6.000 7.350 6.600 8.100 ;
        RECT 4.900 8.300 5.500 9.200 ;
        RECT 7.500 8.450 21.300 9.050 ;
        RECT 20.700 7.550 21.300 9.050 ;
        RECT 4.900 8.600 8.100 9.200 ;
  END 
END dffpr_3

MACRO dffpr_2
  CLASS  CORE ;
  FOREIGN dffpr_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 21.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 15.950 5.950 17.950 6.550 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 5.700 0.000 6.300 2.700 ;
        RECT 0.000 0.000 21.250 2.500 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.100 4.700 1.700 6.250 ;
        RECT 1.100 4.700 2.800 5.400 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 4.450 13.550 5.050 16.250 ;
        RECT 0.000 13.750 21.250 16.250 ;
        RECT 14.450 13.450 15.050 16.250 ;
        RECT 7.950 13.550 8.550 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 12.950 5.950 14.950 6.550 ;
    END
  END qb
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 19.000 8.450 21.000 9.050 ;
    END
  END ck
  PIN rb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.950 7.550 1.550 9.050 ;
        RECT 0.350 8.450 1.550 9.050 ;
    END
  END rb
  OBS 
      LAYER Metal1 ;
        RECT 4.100 5.800 9.800 6.400 ;
        RECT 2.350 6.000 4.700 6.600 ;
        RECT 2.350 6.000 2.950 9.200 ;
        RECT 2.350 8.600 5.250 9.200 ;
        RECT 6.100 8.450 18.500 9.050 ;
        RECT 9.300 8.450 10.000 9.200 ;
        RECT 8.400 7.250 9.100 7.950 ;
        RECT 18.200 7.250 19.800 7.850 ;
        RECT 3.550 7.350 18.800 7.950 ;
        RECT 3.550 7.350 4.150 8.100 ;
        RECT 11.600 3.350 20.050 3.950 ;
  END 
END dffpr_2

MACRO dffpr_1
  CLASS  CORE ;
  FOREIGN dffpr_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 21.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 15.950 5.950 17.950 6.550 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 5.700 0.000 6.300 2.700 ;
        RECT 0.000 0.000 21.250 2.500 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.100 4.700 1.700 6.300 ;
        RECT 1.100 4.700 2.800 5.400 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 4.450 13.550 5.050 16.250 ;
        RECT 0.000 13.750 21.250 16.250 ;
        RECT 7.950 13.550 8.550 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 12.900 5.950 14.900 6.550 ;
    END
  END qb
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 19.000 8.450 21.000 9.050 ;
    END
  END ck
  PIN rb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.950 7.550 1.550 9.050 ;
        RECT 0.350 8.450 1.550 9.050 ;
    END
  END rb
  OBS 
      LAYER Metal1 ;
        RECT 4.100 5.800 9.800 6.400 ;
        RECT 2.350 6.000 4.700 6.600 ;
        RECT 2.350 6.000 2.950 9.200 ;
        RECT 2.350 8.600 5.250 9.200 ;
        RECT 6.100 8.450 18.500 9.050 ;
        RECT 9.300 8.450 10.000 9.200 ;
        RECT 3.550 7.250 19.800 7.850 ;
        RECT 3.550 7.250 4.150 8.100 ;
        RECT 11.600 3.350 20.050 3.950 ;
  END 
END dffpr_1

MACRO dffphc_8
  CLASS  CORE ;
  FOREIGN dffphc_8 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 33.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 28.500 9.700 30.500 10.300 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 33.750 2.500 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.150 8.450 4.150 9.050 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 4.400 13.550 5.000 16.250 ;
        RECT 0.000 13.750 33.750 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 24.850 9.700 26.850 10.300 ;
    END
  END qb
  PIN g
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.400 7.200 5.950 7.800 ;
        RECT 5.350 7.200 5.950 8.350 ;
    END
  END g
  PIN clb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.350 4.700 2.350 5.300 ;
    END
  END clb
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 31.250 4.700 33.250 5.300 ;
    END
  END ck
  OBS 
      LAYER Metal1 ;
        RECT 6.100 4.550 6.700 5.300 ;
        RECT 4.400 4.700 6.700 5.300 ;
        RECT 1.450 5.950 8.400 6.550 ;
        RECT 9.150 6.100 10.100 6.700 ;
        RECT 9.150 6.100 9.750 10.350 ;
        RECT 19.250 5.750 19.850 6.550 ;
        RECT 11.800 5.950 19.850 6.550 ;
        RECT 11.800 5.950 12.400 9.050 ;
        RECT 11.350 8.450 16.750 9.050 ;
        RECT 7.300 4.550 7.900 5.300 ;
        RECT 7.300 4.700 11.200 5.300 ;
        RECT 10.600 4.700 11.200 7.850 ;
        RECT 10.250 7.250 10.850 10.300 ;
        RECT 10.250 9.700 22.950 10.300 ;
        RECT 17.250 4.650 28.450 5.250 ;
        RECT 19.200 7.050 19.800 7.800 ;
        RECT 12.900 7.200 33.150 7.800 ;
  END 
END dffphc_8

MACRO dffphc_6
  CLASS  CORE ;
  FOREIGN dffphc_6 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 32.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 27.000 9.700 29.000 10.300 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 13.900 0.000 14.500 2.800 ;
        RECT 0.000 0.000 32.500 2.500 ;
        RECT 26.300 0.000 26.900 2.800 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.800 8.450 2.950 9.050 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 4.000 13.550 4.600 16.250 ;
        RECT 0.000 13.750 32.500 16.250 ;
        RECT 26.300 13.450 26.900 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 21.600 8.450 23.600 9.050 ;
    END
  END qb
  PIN g
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.850 7.200 5.650 7.800 ;
        RECT 5.050 7.200 5.650 7.950 ;
    END
  END g
  PIN clb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 5.950 2.250 6.550 ;
    END
  END clb
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 30.000 7.200 32.000 7.800 ;
    END
  END ck
  OBS 
      LAYER Metal1 ;
        RECT 5.900 4.550 6.500 5.250 ;
        RECT 4.000 4.650 6.500 5.250 ;
        RECT 1.000 4.700 3.400 5.300 ;
        RECT 2.800 4.700 3.400 6.500 ;
        RECT 2.800 5.900 8.250 6.500 ;
        RECT 7.650 5.900 8.250 10.300 ;
        RECT 1.050 9.700 8.250 10.300 ;
        RECT 9.450 6.100 10.050 10.300 ;
        RECT 10.550 5.950 18.650 6.550 ;
        RECT 10.550 5.950 11.150 8.950 ;
        RECT 10.550 8.350 15.550 8.950 ;
        RECT 13.650 9.500 14.250 10.250 ;
        RECT 13.650 9.650 25.200 10.250 ;
        RECT 7.100 4.550 7.700 5.400 ;
        RECT 7.100 4.800 25.200 5.400 ;
        RECT 20.250 7.100 26.500 7.700 ;
        RECT 20.250 7.100 20.850 9.150 ;
        RECT 16.950 8.550 20.850 9.150 ;
        RECT 19.150 5.950 32.050 6.550 ;
        RECT 19.150 5.950 19.750 7.850 ;
        RECT 11.650 7.250 19.750 7.850 ;
  END 
END dffphc_6

MACRO dffphc_4
  CLASS  CORE ;
  FOREIGN dffphc_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 30.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 24.950 7.200 26.950 7.800 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 6.100 0.000 6.700 2.750 ;
        RECT 0.000 0.000 30.000 2.500 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.200 8.450 4.200 9.050 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 30.000 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 21.250 5.950 23.250 6.550 ;
    END
  END qb
  PIN g
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.950 5.950 1.550 9.050 ;
        RECT 0.950 5.950 1.750 6.550 ;
        RECT 0.550 8.450 1.550 9.050 ;
    END
  END g
  PIN clb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.550 9.700 6.550 10.300 ;
    END
  END clb
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 12.450 5.950 14.450 6.550 ;
    END
  END ck
  OBS 
      LAYER Metal1 ;
        RECT 4.200 6.200 8.250 6.800 ;
        RECT 9.150 5.950 10.350 6.550 ;
        RECT 9.150 5.950 9.750 7.950 ;
        RECT 8.350 7.350 9.750 7.950 ;
        RECT 8.350 7.350 8.950 10.150 ;
        RECT 8.350 9.550 10.350 10.150 ;
        RECT 9.700 8.450 20.100 9.050 ;
        RECT 10.300 7.350 21.450 7.950 ;
        RECT 6.350 7.500 7.800 8.100 ;
        RECT 22.250 8.100 24.050 8.700 ;
        RECT 22.250 8.100 22.850 10.150 ;
        RECT 10.900 9.550 22.850 10.150 ;
        RECT 7.200 7.500 7.800 11.250 ;
        RECT 10.900 9.550 11.500 11.250 ;
        RECT 7.200 10.650 11.500 11.250 ;
  END 
END dffphc_4

MACRO dffphc_3
  CLASS  CORE ;
  FOREIGN dffphc_3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 27.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 23.750 5.950 25.750 6.550 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 6.100 0.000 6.700 2.750 ;
        RECT 0.000 0.000 27.500 2.500 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.850 8.050 3.450 10.300 ;
        RECT 1.850 9.700 3.450 10.300 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 27.500 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 20.750 5.950 22.750 6.550 ;
    END
  END qb
  PIN g
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.350 7.200 0.950 9.550 ;
        RECT 0.350 7.200 1.800 7.800 ;
        RECT 1.200 7.100 1.800 7.800 ;
    END
  END g
  PIN clb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.400 8.450 6.250 10.300 ;
        RECT 4.700 9.700 6.250 10.300 ;
    END
  END clb
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 12.650 5.950 14.650 6.550 ;
    END
  END ck
  OBS 
      LAYER Metal1 ;
        RECT 4.100 6.200 8.300 6.800 ;
        RECT 9.350 6.200 10.250 6.800 ;
        RECT 9.350 6.200 9.950 7.950 ;
        RECT 8.400 7.350 9.950 7.950 ;
        RECT 8.400 7.350 9.000 10.150 ;
        RECT 8.400 9.550 10.250 10.150 ;
        RECT 9.500 8.450 19.800 9.050 ;
        RECT 15.450 6.400 16.050 7.950 ;
        RECT 19.200 7.150 19.800 7.950 ;
        RECT 10.450 7.350 19.800 7.950 ;
        RECT 6.350 7.300 7.900 7.900 ;
        RECT 22.650 7.350 23.250 10.150 ;
        RECT 10.750 9.550 23.250 10.150 ;
        RECT 7.300 7.300 7.900 11.350 ;
        RECT 10.750 9.550 11.350 11.350 ;
        RECT 7.300 10.750 11.350 11.350 ;
  END 
END dffphc_3

MACRO dffphc_2
  CLASS  CORE ;
  FOREIGN dffphc_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 25.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 19.800 8.450 21.800 9.050 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 12.800 0.000 13.400 2.700 ;
        RECT 0.000 0.000 25.000 2.500 ;
        RECT 18.800 0.000 19.400 2.800 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.500 8.450 3.500 9.050 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 12.850 13.550 13.450 16.250 ;
        RECT 0.000 13.750 25.000 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 16.950 8.450 18.950 9.050 ;
    END
  END qb
  PIN g
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.150 7.200 5.300 7.800 ;
        RECT 4.700 8.450 6.500 9.050 ;
        RECT 4.700 7.200 5.300 9.050 ;
    END
  END g
  PIN clb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 3.450 2.250 4.050 ;
    END
  END clb
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 22.750 8.450 24.750 9.050 ;
    END
  END ck
  OBS 
      LAYER Metal1 ;
        RECT 1.000 5.950 7.450 6.550 ;
        RECT 6.850 5.950 7.450 7.250 ;
        RECT 9.700 5.800 10.300 6.550 ;
        RECT 7.950 5.950 10.300 6.550 ;
        RECT 7.950 5.950 8.550 9.200 ;
        RECT 7.950 8.600 10.750 9.200 ;
        RECT 11.000 6.250 15.100 6.850 ;
        RECT 11.000 6.250 11.600 7.650 ;
        RECT 9.050 7.050 11.600 7.650 ;
        RECT 9.050 7.050 9.650 8.100 ;
        RECT 6.400 4.700 16.450 5.300 ;
        RECT 6.400 4.700 7.000 5.450 ;
        RECT 15.850 4.700 16.450 6.750 ;
        RECT 15.850 6.150 19.000 6.750 ;
        RECT 15.800 7.250 24.600 7.850 ;
        RECT 13.200 7.350 16.400 7.950 ;
        RECT 13.200 7.350 13.800 8.750 ;
        RECT 11.250 8.150 13.800 8.750 ;
  END 
END dffphc_2

MACRO dffphc_1
  CLASS  CORE ;
  FOREIGN dffphc_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 25.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 22.750 5.950 24.750 6.550 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 21.400 0.000 22.000 2.700 ;
        RECT 0.000 0.000 25.000 2.500 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.000 8.450 4.000 9.050 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 13.150 13.550 13.750 16.250 ;
        RECT 0.000 13.750 25.000 16.250 ;
        RECT 21.350 13.550 21.950 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 21.000 8.450 23.000 9.050 ;
    END
  END qb
  PIN g
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.050 7.200 6.500 7.800 ;
    END
  END g
  PIN clb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 3.350 1.750 4.150 ;
    END
  END clb
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 13.250 3.450 15.250 4.050 ;
    END
  END ck
  OBS 
      LAYER Metal1 ;
        RECT 6.500 5.200 8.300 5.800 ;
        RECT 6.500 5.200 7.100 6.550 ;
        RECT 1.000 5.950 7.100 6.550 ;
        RECT 9.600 5.800 10.200 7.000 ;
        RECT 7.900 6.400 10.200 7.000 ;
        RECT 7.900 6.400 8.500 9.200 ;
        RECT 7.900 8.600 10.700 9.200 ;
        RECT 10.750 6.250 16.900 6.850 ;
        RECT 10.750 6.250 11.350 8.100 ;
        RECT 9.000 7.500 11.350 8.100 ;
        RECT 16.300 8.450 19.500 9.050 ;
        RECT 11.850 7.350 20.200 7.950 ;
  END 
END dffphc_1

MACRO dffph_8
  CLASS  CORE ;
  FOREIGN dffph_8 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 32.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 27.000 8.450 29.000 9.050 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 3.200 0.000 3.800 2.800 ;
        RECT 0.000 0.000 32.500 2.500 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.350 8.450 2.350 9.050 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 22.750 13.450 23.350 16.250 ;
        RECT 0.000 13.750 32.500 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 23.550 8.450 25.550 9.050 ;
    END
  END qb
  PIN g
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.950 7.200 5.450 7.800 ;
    END
  END g
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 29.950 4.700 31.950 5.300 ;
    END
  END ck
  OBS 
      LAYER Metal1 ;
        RECT 0.450 5.800 7.250 6.400 ;
        RECT 7.800 4.700 9.150 5.300 ;
        RECT 7.800 4.700 8.400 10.150 ;
        RECT 7.800 9.550 9.200 10.150 ;
        RECT 8.900 5.950 16.650 6.550 ;
        RECT 8.900 5.900 9.500 9.050 ;
        RECT 8.900 8.450 14.750 9.050 ;
        RECT 12.650 9.700 21.650 10.300 ;
        RECT 12.650 9.700 13.250 10.350 ;
        RECT 14.500 4.700 27.150 5.300 ;
        RECT 17.050 7.050 17.650 7.800 ;
        RECT 10.000 7.200 31.850 7.800 ;
  END 
END dffph_8

MACRO dffph_6
  CLASS  CORE ;
  FOREIGN dffph_6 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 31.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 25.850 9.700 27.850 10.300 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 3.050 0.000 3.650 2.800 ;
        RECT 0.000 0.000 31.250 2.500 ;
        RECT 25.050 0.000 25.650 2.800 ;
        RECT 18.650 0.000 19.250 2.800 ;
        RECT 11.800 0.000 12.500 2.550 ;
        RECT 7.200 0.000 7.800 2.700 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.400 8.450 2.750 9.050 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 25.050 13.450 25.650 16.250 ;
        RECT 0.000 13.750 31.250 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 20.350 8.450 22.350 9.050 ;
    END
  END qb
  PIN g
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.200 5.950 4.050 6.550 ;
        RECT 3.450 5.950 4.050 9.050 ;
    END
  END g
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 28.750 5.950 30.750 6.550 ;
    END
  END ck
  OBS 
      LAYER Metal1 ;
        RECT 6.000 6.200 6.600 10.300 ;
        RECT 0.450 9.700 7.200 10.300 ;
        RECT 7.750 4.850 8.600 5.450 ;
        RECT 7.750 4.850 8.350 10.300 ;
        RECT 7.750 9.700 8.950 10.300 ;
        RECT 8.850 5.950 17.400 6.550 ;
        RECT 8.850 5.950 9.450 8.950 ;
        RECT 8.850 8.350 13.950 8.950 ;
        RECT 12.450 9.500 13.050 10.250 ;
        RECT 12.450 9.650 23.950 10.250 ;
        RECT 19.000 7.100 25.400 7.700 ;
        RECT 19.000 7.100 19.600 8.950 ;
        RECT 14.800 8.350 19.600 8.950 ;
        RECT 17.900 6.000 27.000 6.600 ;
        RECT 26.400 6.000 27.000 7.800 ;
        RECT 26.400 7.200 30.800 7.800 ;
        RECT 17.900 6.000 18.500 7.850 ;
        RECT 9.950 7.250 18.500 7.850 ;
  END 
END dffph_6

MACRO dffph_4
  CLASS  CORE ;
  FOREIGN dffph_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 28.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 23.700 7.200 25.700 7.800 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 28.750 2.500 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.200 8.450 4.200 9.050 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 28.750 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 20.000 5.950 22.000 6.550 ;
    END
  END qb
  PIN g
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.950 6.750 1.550 9.350 ;
        RECT 0.950 6.750 1.750 7.350 ;
    END
  END g
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 11.200 5.950 13.200 6.550 ;
    END
  END ck
  OBS 
      LAYER Metal1 ;
        RECT 3.700 6.250 7.000 6.850 ;
        RECT 7.550 5.850 8.800 6.450 ;
        RECT 7.550 5.850 8.150 7.950 ;
        RECT 7.050 7.350 7.650 10.150 ;
        RECT 7.050 9.550 8.900 10.150 ;
        RECT 8.150 8.450 18.800 9.050 ;
        RECT 9.050 7.150 9.650 7.950 ;
        RECT 9.050 7.350 20.200 7.950 ;
        RECT 19.300 8.450 22.850 9.050 ;
        RECT 19.300 8.450 19.900 10.150 ;
        RECT 9.650 9.550 19.900 10.150 ;
        RECT 4.900 8.000 5.500 11.250 ;
        RECT 9.650 9.550 10.250 11.250 ;
        RECT 4.900 10.650 10.250 11.250 ;
  END 
END dffph_4

MACRO dffph_3
  CLASS  CORE ;
  FOREIGN dffph_3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 26.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 22.500 5.950 24.500 6.550 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 26.250 2.500 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.700 7.200 4.700 7.800 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 26.250 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 18.800 5.950 20.800 6.550 ;
    END
  END qb
  PIN g
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.950 5.950 1.550 8.950 ;
        RECT 0.950 5.950 1.650 6.550 ;
    END
  END g
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 11.400 5.950 13.400 6.550 ;
    END
  END ck
  OBS 
      LAYER Metal1 ;
        RECT 3.950 5.950 7.200 6.550 ;
        RECT 8.100 5.900 8.950 6.500 ;
        RECT 8.100 5.900 8.700 7.650 ;
        RECT 6.200 7.050 8.700 7.650 ;
        RECT 6.200 7.050 6.800 10.150 ;
        RECT 6.200 9.550 9.000 10.150 ;
        RECT 8.050 8.300 8.650 9.050 ;
        RECT 8.050 8.450 18.500 9.050 ;
        RECT 9.200 7.000 9.800 7.950 ;
        RECT 14.200 6.750 14.800 7.950 ;
        RECT 17.850 7.150 18.500 7.950 ;
        RECT 9.200 7.350 18.500 7.950 ;
        RECT 19.000 7.350 22.050 7.950 ;
        RECT 19.000 7.350 19.600 10.150 ;
        RECT 9.500 9.550 19.600 10.150 ;
        RECT 4.900 8.300 5.500 11.250 ;
        RECT 9.500 9.550 10.100 11.250 ;
        RECT 4.900 10.650 10.100 11.250 ;
  END 
END dffph_3

MACRO dffph_2
  CLASS  CORE ;
  FOREIGN dffph_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 23.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 18.550 8.450 20.550 9.050 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 3.350 0.000 3.950 2.650 ;
        RECT 0.000 0.000 23.750 2.500 ;
        RECT 17.550 0.000 18.150 2.800 ;
        RECT 11.550 0.000 12.150 2.700 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 8.450 2.300 9.050 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 3.450 13.550 4.050 16.250 ;
        RECT 0.000 13.750 23.750 16.250 ;
        RECT 11.600 13.550 12.200 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 15.700 8.450 17.700 9.050 ;
    END
  END qb
  PIN g
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.200 6.450 2.800 7.800 ;
        RECT 3.450 8.450 4.450 9.050 ;
        RECT 3.450 7.200 4.050 9.050 ;
        RECT 2.200 7.200 4.050 7.800 ;
    END
  END g
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 21.500 8.450 23.500 9.050 ;
    END
  END ck
  OBS 
      LAYER Metal1 ;
        RECT 8.450 5.800 9.050 6.550 ;
        RECT 6.250 5.950 9.050 6.550 ;
        RECT 6.250 5.950 6.850 9.200 ;
        RECT 6.250 8.600 9.050 9.200 ;
        RECT 9.750 6.250 13.850 6.850 ;
        RECT 9.750 6.250 10.350 7.650 ;
        RECT 7.350 7.050 10.350 7.650 ;
        RECT 7.350 7.050 7.950 8.100 ;
        RECT 4.950 4.700 15.200 5.300 ;
        RECT 14.600 4.700 15.200 6.750 ;
        RECT 4.950 4.700 5.550 6.600 ;
        RECT 14.600 6.150 17.750 6.750 ;
        RECT 14.550 7.250 23.350 7.850 ;
        RECT 11.950 7.350 15.150 7.950 ;
        RECT 11.950 7.350 12.550 8.750 ;
        RECT 10.000 8.150 12.550 8.750 ;
  END 
END dffph_2

MACRO dffph_1
  CLASS  CORE ;
  FOREIGN dffph_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 23.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 21.500 5.950 23.500 6.550 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 2.950 0.000 3.550 2.700 ;
        RECT 0.000 0.000 23.750 2.500 ;
        RECT 20.150 0.000 20.750 2.700 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.750 8.450 2.750 9.050 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 3.200 13.550 3.800 16.250 ;
        RECT 0.000 13.750 23.750 16.250 ;
        RECT 20.100 13.550 20.700 16.250 ;
        RECT 11.900 13.550 12.500 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 19.650 8.450 21.650 9.050 ;
    END
  END qb
  PIN g
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.750 7.200 5.300 7.800 ;
    END
  END g
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 12.100 3.450 14.100 4.050 ;
    END
  END ck
  OBS 
      LAYER Metal1 ;
        RECT 5.250 5.300 7.000 5.900 ;
        RECT 5.250 5.300 5.850 6.550 ;
        RECT 0.350 5.950 5.850 6.550 ;
        RECT 8.350 5.800 8.950 7.000 ;
        RECT 6.600 6.400 8.950 7.000 ;
        RECT 6.600 6.400 7.200 9.200 ;
        RECT 6.600 8.600 9.400 9.200 ;
        RECT 9.500 6.250 15.650 6.850 ;
        RECT 9.500 6.250 10.100 8.100 ;
        RECT 7.700 7.500 10.100 8.100 ;
        RECT 15.050 8.450 18.250 9.050 ;
        RECT 10.600 7.350 18.950 7.950 ;
  END 
END dffph_1

MACRO dffpc_8
  CLASS  CORE ;
  FOREIGN dffpc_8 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 28.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 23.100 8.450 25.100 9.050 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 28.750 2.500 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.600 8.450 3.700 9.050 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 28.750 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 19.150 8.450 21.150 9.050 ;
    END
  END qb
  PIN clb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.400 7.200 2.400 7.800 ;
    END
  END clb
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 26.050 4.700 28.050 5.300 ;
    END
  END ck
  OBS 
      LAYER Metal1 ;
        RECT 4.200 4.850 5.300 5.450 ;
        RECT 4.200 4.850 4.800 10.300 ;
        RECT 4.200 9.700 5.300 10.300 ;
        RECT 5.300 5.950 14.350 6.550 ;
        RECT 5.300 5.950 5.900 9.050 ;
        RECT 5.300 8.450 10.800 9.050 ;
        RECT 8.900 9.600 9.500 10.300 ;
        RECT 8.900 9.700 17.750 10.300 ;
        RECT 11.250 4.700 23.250 5.300 ;
        RECT 12.950 7.050 13.550 7.800 ;
        RECT 6.400 7.200 27.950 7.800 ;
        RECT 6.400 7.200 7.000 7.850 ;
  END 
END dffpc_8

MACRO dffpc_6
  CLASS  CORE ;
  FOREIGN dffpc_6 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 27.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 22.000 9.700 24.000 10.300 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 21.300 0.000 21.900 2.650 ;
        RECT 0.000 0.000 27.500 2.500 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.350 8.450 2.350 9.050 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 1.000 13.450 1.600 16.250 ;
        RECT 0.000 13.750 27.500 16.250 ;
        RECT 21.300 13.450 21.900 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 16.600 8.450 18.600 9.050 ;
    END
  END qb
  PIN clb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.350 4.700 2.750 5.300 ;
    END
  END clb
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 25.000 5.950 27.000 6.550 ;
    END
  END ck
  OBS 
      LAYER Metal1 ;
        RECT 4.400 5.250 5.000 6.500 ;
        RECT 3.400 5.900 5.000 6.500 ;
        RECT 3.400 5.900 4.000 10.300 ;
        RECT 3.400 9.700 5.200 10.300 ;
        RECT 9.500 8.200 10.100 8.900 ;
        RECT 5.350 8.300 10.100 8.900 ;
        RECT 6.050 5.650 13.650 6.250 ;
        RECT 6.050 5.650 6.650 6.550 ;
        RECT 8.600 9.500 9.200 10.250 ;
        RECT 8.600 9.650 20.200 10.250 ;
        RECT 15.250 7.100 21.300 7.700 ;
        RECT 15.250 7.100 15.850 8.900 ;
        RECT 11.450 8.300 15.850 8.900 ;
        RECT 14.150 6.000 23.250 6.600 ;
        RECT 22.650 6.000 23.250 7.800 ;
        RECT 7.500 7.100 14.750 7.700 ;
        RECT 4.500 7.200 8.100 7.800 ;
        RECT 14.150 6.000 14.750 7.800 ;
        RECT 13.050 7.100 14.750 7.800 ;
        RECT 22.650 7.200 27.050 7.800 ;
  END 
END dffpc_6

MACRO dffpc_4
  CLASS  CORE ;
  FOREIGN dffpc_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 25.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 20.550 7.200 22.550 7.800 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 25.000 2.500 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.950 5.950 2.950 6.550 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 25.000 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 16.750 5.950 18.750 6.550 ;
    END
  END qb
  PIN clb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.350 8.450 2.550 9.050 ;
    END
  END clb
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.450 5.950 9.450 6.550 ;
    END
  END ck
  OBS 
      LAYER Metal1 ;
        RECT 3.600 5.950 5.150 6.550 ;
        RECT 3.600 5.950 4.200 7.850 ;
        RECT 3.250 7.250 3.850 10.550 ;
        RECT 3.250 9.950 5.050 10.550 ;
        RECT 10.650 6.050 15.300 6.650 ;
        RECT 14.700 6.050 15.300 7.100 ;
        RECT 10.650 6.050 11.250 7.950 ;
        RECT 5.200 7.350 11.250 7.950 ;
        RECT 11.850 7.300 12.450 9.050 ;
        RECT 4.400 8.450 16.750 9.050 ;
  END 
END dffpc_4

MACRO dffpc_3
  CLASS  CORE ;
  FOREIGN dffpc_3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 22.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 18.550 5.950 20.550 6.550 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 7.150 0.000 7.750 2.750 ;
        RECT 0.000 0.000 22.500 2.500 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.900 5.950 2.900 6.550 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 22.500 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 15.750 5.950 17.750 6.550 ;
    END
  END qb
  PIN clb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 8.450 2.250 9.050 ;
    END
  END clb
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.950 5.950 9.950 6.550 ;
    END
  END ck
  OBS 
      LAYER Metal1 ;
        RECT 3.500 6.000 5.100 6.600 ;
        RECT 3.500 6.000 4.100 7.950 ;
        RECT 3.000 7.350 3.600 10.350 ;
        RECT 3.000 9.750 5.050 10.350 ;
        RECT 4.350 8.450 15.550 9.050 ;
        RECT 4.350 8.450 4.950 9.250 ;
        RECT 5.000 7.350 15.550 7.950 ;
  END 
END dffpc_3

MACRO dffpc_2
  CLASS  CORE ;
  FOREIGN dffpc_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 20.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 14.800 8.450 16.800 9.050 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 7.800 0.000 8.400 2.700 ;
        RECT 0.000 0.000 20.000 2.500 ;
        RECT 13.800 0.000 14.400 2.800 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.150 4.700 3.500 5.300 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 1.050 13.550 1.650 16.250 ;
        RECT 0.000 13.750 20.000 16.250 ;
        RECT 7.850 13.550 8.450 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 11.950 8.450 13.950 9.050 ;
    END
  END qb
  PIN clb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 8.450 2.250 9.050 ;
    END
  END clb
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 17.750 8.450 19.750 9.050 ;
    END
  END ck
  OBS 
      LAYER Metal1 ;
        RECT 4.700 5.800 5.300 6.550 ;
        RECT 2.900 5.950 5.300 6.550 ;
        RECT 2.900 5.950 3.500 9.200 ;
        RECT 2.900 8.600 5.300 9.200 ;
        RECT 6.000 6.250 10.100 6.850 ;
        RECT 6.000 6.250 6.600 7.650 ;
        RECT 4.000 7.050 6.600 7.650 ;
        RECT 4.000 7.050 4.600 8.100 ;
        RECT 10.800 7.250 19.600 7.850 ;
        RECT 8.200 7.350 11.400 7.950 ;
        RECT 8.200 7.350 8.800 8.750 ;
        RECT 6.250 8.150 8.800 8.750 ;
  END 
END dffpc_2

MACRO dffpc_1
  CLASS  CORE ;
  FOREIGN dffpc_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 18.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 16.500 5.950 18.500 6.550 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 7.350 0.000 7.950 2.700 ;
        RECT 0.000 0.000 18.750 2.500 ;
        RECT 16.050 0.000 16.650 2.700 ;
        RECT 9.950 0.000 10.550 2.700 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.950 4.700 2.950 5.300 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 1.000 13.550 1.600 16.250 ;
        RECT 0.000 13.750 18.750 16.250 ;
        RECT 16.000 13.550 16.600 16.250 ;
        RECT 7.800 13.550 8.400 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 15.250 8.450 17.250 9.050 ;
    END
  END qb
  PIN clb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.950 7.500 1.550 9.050 ;
        RECT 0.350 8.450 1.550 9.050 ;
    END
  END clb
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.300 3.450 9.300 4.050 ;
    END
  END ck
  OBS 
      LAYER Metal1 ;
        RECT 4.250 5.800 4.850 7.000 ;
        RECT 2.500 6.400 4.850 7.000 ;
        RECT 2.500 6.400 3.100 9.200 ;
        RECT 2.500 8.600 5.300 9.200 ;
        RECT 5.500 6.250 11.550 6.850 ;
        RECT 5.500 6.250 6.100 8.100 ;
        RECT 3.600 7.500 6.100 8.100 ;
        RECT 10.950 8.450 14.150 9.050 ;
        RECT 6.600 7.350 14.850 7.950 ;
  END 
END dffpc_1

MACRO dffp_8
  CLASS  CORE ;
  FOREIGN dffp_8 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 26.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 20.600 5.950 22.600 6.550 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 26.250 2.500 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.350 8.450 1.550 9.050 ;
        RECT 0.950 8.450 1.550 10.300 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 16.350 13.450 16.950 16.250 ;
        RECT 0.000 13.750 26.250 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 16.650 8.450 18.650 9.050 ;
    END
  END qb
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 23.550 4.700 25.550 5.300 ;
    END
  END ck
  OBS 
      LAYER Metal1 ;
        RECT 2.550 4.700 3.950 5.300 ;
        RECT 2.550 4.700 3.150 10.300 ;
        RECT 2.550 9.700 3.950 10.300 ;
        RECT 11.200 5.750 11.800 6.400 ;
        RECT 3.650 5.800 11.800 6.400 ;
        RECT 3.650 5.800 5.500 6.550 ;
        RECT 3.650 5.800 4.250 9.000 ;
        RECT 3.650 8.400 9.500 9.000 ;
        RECT 8.900 8.400 9.500 9.050 ;
        RECT 7.600 9.700 15.250 10.300 ;
        RECT 10.000 4.650 20.750 5.250 ;
        RECT 11.200 7.050 11.800 7.850 ;
        RECT 4.750 7.200 25.450 7.850 ;
  END 
END dffp_8

MACRO dffp_6
  CLASS  CORE ;
  FOREIGN dffp_6 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 25.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 19.600 9.700 21.600 10.300 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 18.800 0.000 19.400 2.650 ;
        RECT 0.000 0.000 25.000 2.500 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.350 4.700 1.550 5.300 ;
        RECT 0.950 4.700 1.550 6.300 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 18.800 13.450 19.400 16.250 ;
        RECT 0.000 13.750 25.000 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 14.100 8.450 16.100 9.050 ;
    END
  END qb
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 22.500 5.950 24.500 6.550 ;
    END
  END ck
  OBS 
      LAYER Metal1 ;
        RECT 2.350 4.850 3.800 5.450 ;
        RECT 2.350 4.850 2.950 10.300 ;
        RECT 2.350 9.700 3.550 10.300 ;
        RECT 3.650 5.950 11.150 6.550 ;
        RECT 3.650 5.950 4.250 8.950 ;
        RECT 3.650 8.350 8.950 8.950 ;
        RECT 6.800 9.500 7.400 10.250 ;
        RECT 6.800 9.650 17.700 10.250 ;
        RECT 12.750 7.100 18.800 7.700 ;
        RECT 12.750 7.100 13.350 8.950 ;
        RECT 9.450 8.350 13.350 8.950 ;
        RECT 11.650 5.950 20.750 6.600 ;
        RECT 20.150 5.950 20.750 7.850 ;
        RECT 11.650 5.950 12.250 7.850 ;
        RECT 4.850 7.250 12.250 7.850 ;
        RECT 20.150 7.250 24.550 7.850 ;
  END 
END dffp_6

MACRO dffp_4
  CLASS  CORE ;
  FOREIGN dffp_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 23.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 18.650 7.200 20.650 7.800 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 23.750 2.500 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 4.700 2.250 5.300 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 23.750 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 15.500 5.950 17.500 6.550 ;
    END
  END qb
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.200 5.950 8.200 6.550 ;
    END
  END ck
  OBS 
      LAYER Metal1 ;
        RECT 2.800 5.550 3.900 6.150 ;
        RECT 2.800 5.550 3.400 7.450 ;
        RECT 2.000 6.850 3.400 7.450 ;
        RECT 2.000 6.850 2.600 10.150 ;
        RECT 2.000 9.550 3.800 10.150 ;
        RECT 8.900 6.500 14.400 7.100 ;
        RECT 3.900 6.900 5.300 7.500 ;
        RECT 8.900 6.500 9.500 7.950 ;
        RECT 4.700 7.350 9.500 7.950 ;
        RECT 10.150 7.600 12.600 8.200 ;
        RECT 3.100 8.000 3.700 9.050 ;
        RECT 12.000 7.600 12.600 9.050 ;
        RECT 10.150 7.600 10.750 9.050 ;
        RECT 3.100 8.450 10.750 9.050 ;
        RECT 12.000 8.450 15.500 9.050 ;
  END 
END dffp_4

MACRO dffp_3
  CLASS  CORE ;
  FOREIGN dffp_3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 21.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 17.300 5.950 19.300 6.550 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 5.900 0.000 6.500 2.750 ;
        RECT 0.000 0.000 21.250 2.500 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 4.700 2.250 5.300 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 21.250 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 14.500 5.950 16.500 6.550 ;
    END
  END qb
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.200 5.950 8.200 6.550 ;
    END
  END ck
  OBS 
      LAYER Metal1 ;
        RECT 0.700 5.950 3.800 6.550 ;
        RECT 0.700 5.950 1.300 10.200 ;
        RECT 0.700 9.600 3.800 10.200 ;
        RECT 2.100 8.400 2.700 9.050 ;
        RECT 2.100 8.450 14.500 9.050 ;
        RECT 2.450 7.300 4.300 7.900 ;
        RECT 3.700 7.350 14.500 7.950 ;
  END 
END dffp_3

MACRO dffp_2
  CLASS  CORE ;
  FOREIGN dffp_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 18.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 13.550 8.450 15.550 9.050 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 6.550 0.000 7.150 2.700 ;
        RECT 0.000 0.000 18.750 2.500 ;
        RECT 12.550 0.000 13.150 2.800 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 3.450 2.250 4.050 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 6.600 13.550 7.200 16.250 ;
        RECT 0.000 13.750 18.750 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 10.700 8.450 12.700 9.050 ;
    END
  END qb
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 16.450 8.450 18.450 9.050 ;
    END
  END ck
  OBS 
      LAYER Metal1 ;
        RECT 3.450 5.800 4.050 6.550 ;
        RECT 1.250 5.950 4.050 6.550 ;
        RECT 1.250 5.950 1.850 9.200 ;
        RECT 1.250 8.600 4.050 9.200 ;
        RECT 4.750 6.250 8.850 6.850 ;
        RECT 4.750 6.250 5.350 7.650 ;
        RECT 2.350 7.050 5.350 7.650 ;
        RECT 2.350 7.050 2.950 8.100 ;
        RECT 9.550 7.250 18.350 7.850 ;
        RECT 6.950 7.350 10.150 7.950 ;
        RECT 6.950 7.350 7.550 8.750 ;
        RECT 5.000 8.150 7.550 8.750 ;
  END 
END dffp_2

MACRO dffp_1
  CLASS  CORE ;
  FOREIGN dffp_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 17.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 15.250 5.950 17.250 6.550 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 6.100 0.000 6.700 2.700 ;
        RECT 0.000 0.000 17.500 2.500 ;
        RECT 14.800 0.000 15.400 2.700 ;
        RECT 8.700 0.000 9.300 2.700 ;
    END
  END vss!
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 3.450 2.250 4.050 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 6.550 13.550 7.150 16.250 ;
        RECT 0.000 13.750 17.500 16.250 ;
        RECT 14.750 13.550 15.350 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 14.000 8.450 16.000 9.050 ;
    END
  END qb
  PIN ck
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.550 3.450 8.550 4.050 ;
    END
  END ck
  OBS 
      LAYER Metal1 ;
        RECT 3.000 5.800 3.600 6.550 ;
        RECT 1.250 5.950 3.600 6.550 ;
        RECT 1.250 5.950 1.850 9.200 ;
        RECT 1.250 8.600 4.050 9.200 ;
        RECT 4.250 6.250 10.300 6.850 ;
        RECT 4.250 6.250 4.850 8.100 ;
        RECT 2.350 7.500 4.850 8.100 ;
        RECT 9.700 8.450 12.900 9.050 ;
        RECT 5.350 7.350 13.600 7.950 ;
  END 
END dffp_1

MACRO dffnr_8
  CLASS  CORE ;
  FOREIGN dffnr_8 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 28.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 17.200 9.700 21.200 10.300 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 18.900 0.000 19.500 2.800 ;
        RECT 0.000 0.000 28.750 2.500 ;
    END
  END vss!
  PIN ckb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 26.100 4.700 28.100 5.300 ;
    END
  END ckb
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.950 5.950 2.950 6.550 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 7.250 13.450 7.850 16.250 ;
        RECT 0.000 13.750 28.750 16.250 ;
        RECT 25.700 13.450 26.300 16.250 ;
        RECT 18.900 13.450 19.500 16.250 ;
        RECT 14.200 13.450 14.800 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 23.150 8.450 25.650 9.050 ;
    END
  END qb
  PIN rb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.300 8.450 2.300 9.050 ;
    END
  END rb
  OBS 
      LAYER Metal1 ;
        RECT 3.450 5.150 5.000 5.750 ;
        RECT 3.450 5.150 4.050 10.450 ;
        RECT 3.450 9.850 5.400 10.450 ;
        RECT 6.000 7.350 10.500 7.950 ;
        RECT 7.750 4.550 15.400 5.150 ;
        RECT 7.750 4.550 8.350 5.750 ;
        RECT 14.800 4.550 15.400 6.600 ;
        RECT 8.650 9.550 9.250 10.450 ;
        RECT 8.650 9.850 16.500 10.450 ;
        RECT 11.200 6.750 11.850 7.350 ;
        RECT 11.250 6.750 11.850 9.350 ;
        RECT 16.050 8.450 19.850 9.050 ;
        RECT 11.250 8.750 16.650 9.350 ;
        RECT 17.600 5.300 23.300 5.900 ;
        RECT 8.850 5.650 13.450 6.250 ;
        RECT 4.550 6.250 9.450 6.850 ;
        RECT 12.850 5.650 13.450 7.800 ;
        RECT 12.850 7.200 28.000 7.800 ;
        RECT 4.550 6.250 5.150 9.050 ;
        RECT 4.550 8.450 10.550 9.050 ;
        RECT 9.950 8.450 10.550 9.200 ;
  END 
END dffnr_8

MACRO dffnr_6
  CLASS  CORE ;
  FOREIGN dffnr_6 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 26.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 20.850 9.700 22.850 10.300 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 20.150 0.000 20.750 2.800 ;
        RECT 0.000 0.000 26.250 2.500 ;
        RECT 23.550 0.000 24.150 2.800 ;
    END
  END vss!
  PIN ckb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 23.750 4.700 25.750 5.300 ;
    END
  END ckb
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.500 5.950 2.900 6.550 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 7.200 13.450 7.800 16.250 ;
        RECT 0.000 13.750 26.250 16.250 ;
        RECT 20.100 13.450 20.700 16.250 ;
        RECT 17.100 13.450 17.700 16.250 ;
        RECT 13.700 13.450 14.300 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 15.850 5.950 18.150 6.550 ;
    END
  END qb
  PIN rb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.350 8.450 2.350 9.050 ;
    END
  END rb
  OBS 
      LAYER Metal1 ;
        RECT 4.500 5.650 5.100 7.300 ;
        RECT 4.600 6.700 5.200 9.350 ;
        RECT 5.900 7.350 10.000 7.950 ;
        RECT 5.900 7.350 6.500 8.600 ;
        RECT 7.350 4.550 14.850 5.150 ;
        RECT 7.350 4.550 7.950 5.750 ;
        RECT 14.250 4.550 14.850 5.950 ;
        RECT 8.100 9.550 8.700 10.450 ;
        RECT 8.100 9.850 19.000 10.450 ;
        RECT 10.700 6.750 11.300 9.050 ;
        RECT 10.700 8.450 23.750 9.050 ;
        RECT 3.400 4.550 6.600 5.150 ;
        RECT 6.000 4.550 6.600 6.850 ;
        RECT 8.600 5.650 12.400 6.250 ;
        RECT 6.000 6.250 9.200 6.850 ;
        RECT 11.800 6.250 13.850 6.850 ;
        RECT 13.250 6.250 13.850 7.950 ;
        RECT 3.400 4.550 4.000 10.450 ;
        RECT 13.250 7.350 25.850 7.950 ;
        RECT 7.000 8.450 10.000 9.050 ;
        RECT 9.400 8.450 10.000 9.250 ;
        RECT 3.400 7.850 4.100 10.450 ;
        RECT 7.000 8.450 7.600 10.450 ;
        RECT 3.400 9.850 7.600 10.450 ;
  END 
END dffnr_6

MACRO dffnr_4
  CLASS  CORE ;
  FOREIGN dffnr_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 22.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 16.550 9.700 18.550 10.300 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 22.500 2.500 ;
    END
  END vss!
  PIN ckb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 21.550 6.850 22.150 10.300 ;
        RECT 20.750 9.700 22.150 10.300 ;
    END
  END ckb
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.100 5.950 3.100 6.550 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 22.500 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 13.050 9.700 15.050 10.300 ;
    END
  END qb
  PIN rb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 8.450 2.250 9.050 ;
    END
  END rb
  OBS 
      LAYER Metal1 ;
        RECT 4.000 6.100 10.500 6.700 ;
        RECT 4.000 6.100 4.600 7.800 ;
        RECT 3.300 7.200 4.600 7.800 ;
        RECT 3.300 7.200 3.900 10.300 ;
        RECT 3.300 9.700 5.850 10.300 ;
        RECT 4.400 8.300 5.000 9.050 ;
        RECT 19.300 6.400 19.900 9.050 ;
        RECT 4.400 8.450 19.900 9.050 ;
        RECT 17.900 4.700 21.300 5.300 ;
        RECT 12.600 6.200 13.200 7.950 ;
        RECT 17.900 4.700 18.500 7.950 ;
        RECT 5.600 7.350 18.500 7.950 ;
        RECT 20.400 4.700 21.000 8.600 ;
  END 
END dffnr_4

MACRO dffnr_3
  CLASS  CORE ;
  FOREIGN dffnr_3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 22.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 16.300 5.950 18.300 6.550 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 22.500 2.500 ;
    END
  END vss!
  PIN ckb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 21.550 5.000 22.150 6.550 ;
        RECT 20.250 5.950 22.150 6.550 ;
    END
  END ckb
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.100 5.950 3.400 6.550 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 22.500 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 13.450 9.700 15.450 10.300 ;
    END
  END qb
  PIN rb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 8.450 2.250 9.050 ;
    END
  END rb
  OBS 
      LAYER Metal1 ;
        RECT 4.400 6.100 10.350 6.700 ;
        RECT 4.400 6.100 5.000 7.800 ;
        RECT 3.500 7.200 5.000 7.800 ;
        RECT 3.500 7.200 4.100 10.300 ;
        RECT 3.500 9.700 5.100 10.300 ;
        RECT 4.900 8.300 5.500 9.200 ;
        RECT 7.500 8.450 19.750 9.050 ;
        RECT 4.900 8.600 8.100 9.200 ;
        RECT 12.550 6.350 13.150 7.950 ;
        RECT 6.000 7.350 21.300 7.950 ;
        RECT 6.000 7.350 6.600 8.100 ;
  END 
END dffnr_3

MACRO dffnr_2
  CLASS  CORE ;
  FOREIGN dffnr_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 21.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 15.950 5.950 16.650 9.300 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 14.500 0.000 15.100 2.650 ;
        RECT 0.000 0.000 21.250 2.500 ;
    END
  END vss!
  PIN ckb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 19.700 7.650 20.300 9.050 ;
        RECT 19.700 8.450 21.000 9.050 ;
    END
  END ckb
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.150 5.950 3.450 6.550 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 8.250 13.550 8.850 16.250 ;
        RECT 0.000 13.750 21.250 16.250 ;
        RECT 14.750 13.450 15.350 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 13.050 5.950 13.650 9.300 ;
        RECT 13.050 5.950 14.050 6.550 ;
    END
  END qb
  PIN rb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 8.450 2.250 9.050 ;
    END
  END rb
  OBS 
      LAYER Metal1 ;
        RECT 6.300 7.350 10.300 7.950 ;
        RECT 6.300 7.350 6.950 8.100 ;
        RECT 4.500 6.200 10.300 6.800 ;
        RECT 4.500 6.200 5.100 7.800 ;
        RECT 3.550 7.200 5.100 7.800 ;
        RECT 3.550 7.200 4.150 10.450 ;
        RECT 3.550 9.850 5.300 10.450 ;
        RECT 10.800 4.750 11.450 9.300 ;
        RECT 4.650 8.650 9.450 9.250 ;
        RECT 8.850 8.450 9.450 10.400 ;
        RECT 11.950 8.400 12.550 10.400 ;
        RECT 17.150 7.900 17.750 10.400 ;
        RECT 8.850 9.800 17.750 10.400 ;
        RECT 11.950 4.750 19.900 5.350 ;
        RECT 11.950 4.750 12.550 6.800 ;
        RECT 19.300 4.750 19.900 7.100 ;
        RECT 18.400 6.500 19.900 7.100 ;
        RECT 18.400 6.500 19.000 10.400 ;
        RECT 18.400 9.800 19.900 10.400 ;
  END 
END dffnr_2

MACRO dffnr_1
  CLASS  CORE ;
  FOREIGN dffnr_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 21.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 15.750 5.950 17.750 6.550 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 14.500 0.000 15.100 2.650 ;
        RECT 0.000 0.000 21.250 2.500 ;
    END
  END vss!
  PIN ckb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 19.600 8.450 21.000 9.050 ;
        RECT 20.400 8.450 21.000 10.150 ;
    END
  END ckb
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.100 5.950 3.100 6.550 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 8.250 13.550 8.850 16.250 ;
        RECT 0.000 13.750 21.250 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 13.050 5.950 15.050 6.550 ;
    END
  END qb
  PIN rb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 8.450 2.250 9.050 ;
    END
  END rb
  OBS 
      LAYER Metal1 ;
        RECT 3.900 6.100 10.200 6.700 ;
        RECT 3.900 6.100 4.500 10.450 ;
        RECT 3.900 9.850 5.100 10.450 ;
        RECT 9.750 7.200 10.350 7.950 ;
        RECT 5.450 7.350 10.350 7.950 ;
        RECT 5.450 7.350 7.000 8.050 ;
        RECT 10.850 5.900 11.500 6.500 ;
        RECT 10.850 5.900 11.450 8.900 ;
        RECT 11.950 8.450 18.000 9.050 ;
        RECT 5.000 8.550 9.450 9.150 ;
        RECT 8.850 8.550 9.450 10.000 ;
        RECT 11.950 8.450 12.550 10.000 ;
        RECT 8.850 9.400 12.550 10.000 ;
        RECT 11.950 7.000 12.550 7.800 ;
        RECT 19.200 6.950 19.800 7.800 ;
        RECT 11.950 7.200 19.800 7.800 ;
        RECT 18.500 7.200 19.100 10.300 ;
        RECT 18.500 9.700 19.800 10.300 ;
  END 
END dffnr_1

MACRO dffnh_8
  CLASS  CORE ;
  FOREIGN dffnh_8 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 31.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 25.750 8.450 27.750 9.050 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 3.050 0.000 3.650 2.800 ;
        RECT 0.000 0.000 31.250 2.500 ;
    END
  END vss!
  PIN ckb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 28.700 4.700 30.700 5.300 ;
    END
  END ckb
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 8.450 2.250 9.050 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 21.500 13.450 22.100 16.250 ;
        RECT 0.000 13.750 31.250 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 22.300 8.450 24.300 9.050 ;
    END
  END qb
  PIN g
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.300 6.400 2.900 7.800 ;
        RECT 3.450 8.500 4.100 9.100 ;
        RECT 3.450 7.100 4.050 9.100 ;
        RECT 2.300 7.100 4.050 7.800 ;
    END
  END g
  OBS 
      LAYER Metal1 ;
        RECT 0.350 5.000 6.250 5.600 ;
        RECT 0.350 5.000 0.950 6.400 ;
        RECT 8.050 6.100 8.650 9.350 ;
        RECT 8.050 8.750 9.150 9.350 ;
        RECT 14.250 7.050 14.850 7.800 ;
        RECT 11.000 7.200 14.850 7.800 ;
        RECT 4.800 7.200 5.400 10.450 ;
        RECT 13.500 9.600 14.100 10.450 ;
        RECT 4.800 9.850 20.400 10.450 ;
        RECT 18.200 5.700 26.050 6.300 ;
        RECT 15.150 5.900 16.000 6.500 ;
        RECT 15.400 5.900 16.000 9.050 ;
        RECT 18.200 5.700 18.800 9.050 ;
        RECT 15.400 8.450 18.800 9.050 ;
        RECT 9.350 4.550 27.300 5.150 ;
        RECT 26.700 4.550 27.300 6.550 ;
        RECT 16.650 4.550 17.250 6.550 ;
        RECT 26.700 5.950 30.600 6.550 ;
        RECT 9.350 4.550 9.950 6.850 ;
        RECT 9.850 6.250 10.450 9.050 ;
  END 
END dffnh_8

MACRO dffnh_6
  CLASS  CORE ;
  FOREIGN dffnh_6 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 30.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 24.600 9.700 26.600 10.300 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 3.050 0.000 3.650 2.800 ;
        RECT 0.000 0.000 30.000 2.500 ;
        RECT 23.800 0.000 24.400 2.800 ;
        RECT 17.400 0.000 18.000 2.700 ;
        RECT 6.700 0.000 7.300 2.700 ;
    END
  END vss!
  PIN ckb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 27.500 5.950 29.500 6.550 ;
    END
  END ckb
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 8.450 2.250 9.050 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 23.800 13.550 24.400 16.250 ;
        RECT 0.000 13.750 30.000 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 19.100 8.450 21.100 9.050 ;
    END
  END qb
  PIN g
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.300 5.950 4.750 6.550 ;
        RECT 4.150 5.950 4.750 9.150 ;
    END
  END g
  OBS 
      LAYER Metal1 ;
        RECT 1.200 4.750 6.500 5.350 ;
        RECT 1.200 4.750 1.800 7.750 ;
        RECT 1.200 7.150 3.350 7.750 ;
        RECT 2.750 7.150 3.350 10.300 ;
        RECT 0.450 9.700 7.100 10.300 ;
        RECT 13.350 6.800 13.950 7.800 ;
        RECT 7.100 7.200 13.950 7.800 ;
        RECT 9.850 7.200 10.450 8.350 ;
        RECT 12.050 9.850 22.700 10.450 ;
        RECT 17.750 7.100 24.000 7.700 ;
        RECT 14.450 5.700 15.050 9.350 ;
        RECT 17.750 7.100 18.350 9.350 ;
        RECT 14.450 8.750 18.350 9.350 ;
        RECT 9.550 4.600 16.150 5.200 ;
        RECT 15.550 4.600 16.150 6.550 ;
        RECT 9.550 4.600 10.150 6.550 ;
        RECT 6.000 5.950 10.150 6.550 ;
        RECT 15.550 5.950 25.750 6.550 ;
        RECT 25.150 5.950 25.750 7.800 ;
        RECT 25.150 7.200 29.550 7.800 ;
        RECT 6.000 5.950 6.600 9.200 ;
        RECT 10.950 8.300 13.950 8.900 ;
        RECT 6.000 8.600 8.200 9.200 ;
        RECT 7.600 8.600 8.200 10.300 ;
        RECT 10.950 8.300 11.550 10.300 ;
        RECT 7.600 9.700 11.550 10.300 ;
  END 
END dffnh_6

MACRO dffnh_4
  CLASS  CORE ;
  FOREIGN dffnh_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 28.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 23.700 7.200 25.700 7.800 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 28.750 2.500 ;
    END
  END vss!
  PIN ckb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 11.200 5.950 13.200 6.550 ;
    END
  END ckb
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.250 7.200 4.250 7.800 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 28.750 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 20.000 5.950 22.000 6.550 ;
    END
  END qb
  PIN g
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.950 6.750 1.550 9.350 ;
        RECT 0.950 6.750 1.600 7.350 ;
        RECT 0.700 8.750 1.550 9.350 ;
    END
  END g
  OBS 
      LAYER Metal1 ;
        RECT 3.750 5.850 7.000 6.450 ;
        RECT 7.500 6.250 8.800 6.850 ;
        RECT 7.500 6.250 8.100 7.950 ;
        RECT 6.200 7.350 8.100 7.950 ;
        RECT 6.200 7.350 6.800 10.150 ;
        RECT 6.200 9.550 8.800 10.150 ;
        RECT 15.000 6.600 15.700 7.950 ;
        RECT 9.200 7.350 18.550 7.950 ;
        RECT 8.050 8.450 19.900 9.050 ;
        RECT 22.200 8.100 22.800 10.150 ;
        RECT 10.000 9.550 22.800 10.150 ;
        RECT 4.800 8.050 5.400 11.250 ;
        RECT 10.000 9.550 10.600 11.250 ;
        RECT 4.800 10.650 10.600 11.250 ;
  END 
END dffnh_4

MACRO dffnh_3
  CLASS  CORE ;
  FOREIGN dffnh_3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 26.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 22.500 5.950 24.500 6.550 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 26.250 2.500 ;
    END
  END vss!
  PIN ckb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 11.400 5.950 13.400 6.550 ;
    END
  END ckb
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.200 7.200 4.200 7.800 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 26.250 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 19.300 5.950 21.300 6.550 ;
    END
  END qb
  PIN g
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.950 5.950 1.550 9.050 ;
        RECT 0.950 5.950 1.650 6.550 ;
        RECT 0.900 8.450 1.550 9.050 ;
    END
  END g
  OBS 
      LAYER Metal1 ;
        RECT 3.950 5.850 7.200 6.450 ;
        RECT 7.700 6.250 9.050 6.850 ;
        RECT 7.700 6.250 8.300 7.950 ;
        RECT 7.150 7.350 7.750 10.150 ;
        RECT 7.150 9.550 9.000 10.150 ;
        RECT 15.250 6.200 15.850 7.950 ;
        RECT 18.650 7.150 19.250 7.950 ;
        RECT 9.250 7.350 19.250 7.950 ;
        RECT 8.250 8.450 19.700 9.050 ;
        RECT 21.400 7.350 22.000 10.150 ;
        RECT 9.500 9.550 22.000 10.150 ;
        RECT 4.900 7.600 5.500 11.250 ;
        RECT 9.500 9.550 10.100 11.250 ;
        RECT 4.900 10.650 10.100 11.250 ;
  END 
END dffnh_3

MACRO dffnh_2
  CLASS  CORE ;
  FOREIGN dffnh_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 23.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 18.600 8.450 20.600 9.050 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 3.100 0.000 3.700 2.650 ;
        RECT 0.000 0.000 23.750 2.500 ;
        RECT 11.550 0.000 12.150 2.700 ;
    END
  END vss!
  PIN ckb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 21.100 8.450 23.100 9.050 ;
    END
  END ckb
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 7.200 2.250 7.800 ;
        RECT 1.650 7.200 2.250 8.250 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 3.450 13.550 4.100 16.250 ;
        RECT 0.000 13.750 23.750 16.250 ;
        RECT 17.950 13.500 18.650 16.250 ;
        RECT 11.900 13.550 12.500 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 16.100 8.450 18.100 9.050 ;
    END
  END qb
  PIN g
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.850 6.450 3.450 7.800 ;
        RECT 3.800 7.200 4.400 9.050 ;
        RECT 2.850 7.200 4.400 7.800 ;
    END
  END g
  OBS 
      LAYER Metal1 ;
        RECT 0.350 9.550 6.800 10.150 ;
        RECT 4.950 5.150 9.100 5.750 ;
        RECT 4.950 5.150 5.550 9.050 ;
        RECT 4.950 8.450 7.900 9.050 ;
        RECT 7.300 8.450 7.900 10.250 ;
        RECT 7.300 9.650 8.900 10.250 ;
        RECT 11.250 6.600 14.250 7.200 ;
        RECT 11.250 6.600 11.850 7.950 ;
        RECT 7.150 7.350 11.850 7.950 ;
        RECT 10.050 5.500 18.050 6.100 ;
        RECT 17.450 5.500 18.050 6.750 ;
        RECT 10.050 5.500 10.650 6.850 ;
        RECT 6.050 6.250 10.650 6.850 ;
        RECT 6.050 6.250 6.650 7.950 ;
        RECT 15.000 7.250 23.400 7.850 ;
        RECT 12.350 7.700 15.600 8.300 ;
        RECT 15.000 7.250 15.600 8.700 ;
        RECT 12.350 7.700 12.950 9.050 ;
        RECT 8.400 8.450 12.950 9.050 ;
        RECT 8.400 8.450 9.000 9.150 ;
  END 
END dffnh_2

MACRO dffnh_1
  CLASS  CORE ;
  FOREIGN dffnh_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 23.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 21.500 5.950 23.500 6.550 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 2.450 0.000 3.050 2.700 ;
        RECT 0.000 0.000 23.750 2.500 ;
        RECT 20.200 0.000 20.800 2.700 ;
    END
  END vss!
  PIN ckb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 10.450 3.450 14.050 4.050 ;
    END
  END ckb
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 7.200 2.250 7.800 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 1.000 13.550 1.600 16.250 ;
        RECT 0.000 13.750 23.750 16.250 ;
        RECT 20.250 13.550 20.850 16.250 ;
        RECT 12.200 13.550 12.800 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 20.350 6.750 20.950 9.050 ;
        RECT 20.100 8.450 21.700 9.050 ;
    END
  END qb
  PIN g
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.400 7.200 5.400 7.800 ;
    END
  END g
  OBS 
      LAYER Metal1 ;
        RECT 1.650 8.450 7.000 9.050 ;
        RECT 8.200 3.400 8.800 4.050 ;
        RECT 3.600 3.450 8.800 4.050 ;
        RECT 7.500 5.850 9.200 6.450 ;
        RECT 7.500 5.850 8.100 10.150 ;
        RECT 7.500 9.550 9.200 10.150 ;
        RECT 9.550 8.250 10.150 9.050 ;
        RECT 14.050 8.400 18.650 9.000 ;
        RECT 17.850 8.250 18.650 9.000 ;
        RECT 9.550 8.450 14.650 9.050 ;
        RECT 8.600 6.950 11.250 7.550 ;
        RECT 15.350 7.150 19.000 7.750 ;
        RECT 10.650 7.300 15.950 7.900 ;
        RECT 10.650 6.950 11.250 7.950 ;
  END 
END dffnh_1

MACRO dffn_8
  CLASS  CORE ;
  FOREIGN dffn_8 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 26.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 20.950 9.700 22.950 10.300 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 6.250 0.000 6.850 2.800 ;
        RECT 0.000 0.000 26.250 2.500 ;
    END
  END vss!
  PIN ckb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 23.550 4.700 25.550 5.300 ;
    END
  END ckb
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.350 8.450 1.550 9.050 ;
        RECT 0.950 8.450 1.550 9.850 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 16.350 13.450 16.950 16.250 ;
        RECT 0.000 13.750 26.250 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 16.650 9.700 18.650 10.300 ;
    END
  END qb
  OBS 
      LAYER Metal1 ;
        RECT 2.550 4.850 3.950 5.450 ;
        RECT 2.550 4.850 3.150 10.350 ;
        RECT 2.550 9.750 3.950 10.350 ;
        RECT 4.800 7.350 11.400 7.950 ;
        RECT 6.700 9.700 15.250 10.300 ;
        RECT 9.800 4.700 20.750 5.300 ;
        RECT 3.700 6.050 11.550 6.650 ;
        RECT 3.700 6.050 4.300 9.050 ;
        RECT 3.700 8.450 25.450 9.050 ;
  END 
END dffn_8

MACRO dffn_6
  CLASS  CORE ;
  FOREIGN dffn_6 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 25.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 19.600 9.700 21.600 10.300 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 18.800 0.000 19.400 2.650 ;
        RECT 0.000 0.000 25.000 2.500 ;
    END
  END vss!
  PIN ckb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 22.650 5.950 24.650 6.550 ;
    END
  END ckb
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 4.700 1.550 5.300 ;
        RECT 0.950 4.700 1.550 6.300 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 18.800 13.450 19.400 16.250 ;
        RECT 0.000 13.750 25.000 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 14.100 9.700 16.100 10.300 ;
    END
  END qb
  OBS 
      LAYER Metal1 ;
        RECT 2.400 4.800 3.750 5.400 ;
        RECT 2.400 4.800 3.000 10.300 ;
        RECT 2.400 9.700 3.800 10.300 ;
        RECT 10.550 7.050 11.150 7.800 ;
        RECT 4.700 7.200 11.150 7.800 ;
        RECT 12.900 8.400 17.700 9.000 ;
        RECT 6.600 9.400 7.200 10.300 ;
        RECT 12.900 8.400 13.500 10.300 ;
        RECT 6.600 9.700 13.500 10.300 ;
        RECT 11.700 7.100 19.000 7.700 ;
        RECT 11.700 7.100 12.300 8.900 ;
        RECT 9.450 8.300 12.300 8.900 ;
        RECT 10.700 5.750 20.750 6.350 ;
        RECT 3.600 5.900 11.300 6.500 ;
        RECT 20.150 5.750 20.750 7.800 ;
        RECT 20.150 7.200 24.550 7.800 ;
        RECT 3.600 5.900 4.200 8.900 ;
        RECT 3.600 8.300 8.750 8.900 ;
        RECT 8.150 8.300 8.750 9.200 ;
  END 
END dffn_6

MACRO dffn_4
  CLASS  CORE ;
  FOREIGN dffn_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 23.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 18.650 7.200 20.650 7.800 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 23.750 2.500 ;
    END
  END vss!
  PIN ckb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.200 5.950 7.800 6.950 ;
        RECT 6.700 5.950 8.450 6.550 ;
    END
  END ckb
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 4.700 2.250 5.300 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 23.750 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 15.500 5.950 17.500 6.550 ;
    END
  END qb
  OBS 
      LAYER Metal1 ;
        RECT 2.000 6.250 3.850 6.850 ;
        RECT 2.000 6.250 2.600 10.150 ;
        RECT 2.000 9.550 3.850 10.150 ;
        RECT 3.100 8.450 5.600 9.050 ;
        RECT 13.350 8.450 14.400 9.050 ;
        RECT 5.000 8.450 5.600 9.700 ;
        RECT 13.350 8.450 13.950 9.700 ;
        RECT 5.000 9.100 13.950 9.700 ;
        RECT 4.000 7.350 6.700 7.950 ;
        RECT 12.000 7.350 14.700 7.950 ;
        RECT 6.100 7.750 12.600 8.350 ;
  END 
END dffn_4

MACRO dffn_3
  CLASS  CORE ;
  FOREIGN dffn_3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 21.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 18.000 5.950 20.000 6.550 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 21.250 2.500 ;
    END
  END vss!
  PIN ckb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.800 5.950 7.800 6.550 ;
    END
  END ckb
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 4.700 2.250 5.300 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 21.250 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 14.700 5.950 16.700 6.550 ;
    END
  END qb
  OBS 
      LAYER Metal1 ;
        RECT 0.900 6.250 3.850 6.850 ;
        RECT 0.900 6.250 1.500 10.150 ;
        RECT 0.900 9.550 3.800 10.150 ;
        RECT 3.050 8.450 13.250 9.050 ;
        RECT 3.950 7.350 14.100 7.950 ;
  END 
END dffn_3

MACRO dffn_2
  CLASS  CORE ;
  FOREIGN dffn_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 18.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 14.050 8.450 16.050 9.050 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 6.600 0.000 7.200 2.700 ;
        RECT 0.000 0.000 18.750 2.500 ;
        RECT 12.600 0.000 13.200 2.800 ;
    END
  END vss!
  PIN ckb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 16.600 8.000 17.200 9.050 ;
        RECT 16.600 8.450 18.150 9.050 ;
    END
  END ckb
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 3.450 2.250 4.050 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 6.900 13.550 7.500 16.250 ;
        RECT 0.000 13.750 18.750 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 11.150 8.450 13.500 9.050 ;
    END
  END qb
  OBS 
      LAYER Metal1 ;
        RECT 1.050 5.950 3.850 6.550 ;
        RECT 1.050 5.950 1.650 10.300 ;
        RECT 1.050 9.700 5.100 10.300 ;
        RECT 5.300 6.900 9.200 7.500 ;
        RECT 2.150 7.350 5.950 7.950 ;
        RECT 9.800 6.850 18.400 7.450 ;
        RECT 6.800 8.000 10.500 8.600 ;
        RECT 9.800 6.850 10.500 8.600 ;
        RECT 3.200 8.450 7.400 9.050 ;
  END 
END dffn_2

MACRO dffn_1
  CLASS  CORE ;
  FOREIGN dffn_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 17.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 15.250 5.950 17.250 6.550 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 14.800 0.000 15.400 2.700 ;
        RECT 0.000 0.000 17.500 2.500 ;
    END
  END vss!
  PIN ckb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.600 3.450 8.450 4.050 ;
    END
  END ckb
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.350 3.000 0.950 4.050 ;
        RECT 0.350 3.450 2.050 4.050 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 6.800 13.550 7.400 16.250 ;
        RECT 0.000 13.750 17.500 16.250 ;
        RECT 14.750 13.550 15.350 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 14.000 8.450 16.000 9.050 ;
    END
  END qb
  OBS 
      LAYER Metal1 ;
        RECT 1.000 5.800 3.800 6.400 ;
        RECT 1.000 5.800 1.600 10.150 ;
        RECT 1.000 9.550 3.800 10.150 ;
        RECT 4.100 8.250 4.700 9.050 ;
        RECT 4.100 8.450 12.750 9.050 ;
        RECT 12.050 8.550 13.200 9.200 ;
        RECT 2.100 7.150 5.800 7.750 ;
        RECT 5.200 7.350 13.500 7.950 ;
  END 
END dffn_1

MACRO deche4_8
  CLASS  CORE ;
  FOREIGN deche4_8 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 41.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 20.300 0.000 20.900 2.700 ;
        RECT 0.000 0.000 41.250 2.500 ;
    END
  END vss!
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 2.150 13.550 2.750 16.250 ;
        RECT 0.000 13.750 41.250 16.250 ;
        RECT 38.500 13.550 39.100 16.250 ;
        RECT 35.100 13.550 35.700 16.250 ;
        RECT 31.700 13.550 32.300 16.250 ;
        RECT 28.300 13.550 28.900 16.250 ;
        RECT 24.900 13.550 25.500 16.250 ;
        RECT 15.750 13.550 16.350 16.250 ;
        RECT 12.350 13.550 12.950 16.250 ;
        RECT 8.950 13.550 9.550 16.250 ;
        RECT 5.550 13.550 6.150 16.250 ;
    END
  END vdd!
  PIN sl0
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 19.500 4.700 21.200 5.400 ;
        RECT 20.600 4.700 21.200 5.600 ;
    END
  END sl0
  PIN en
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.500 5.950 19.300 6.550 ;
        RECT 21.950 5.950 39.500 6.550 ;
        RECT 18.700 6.100 22.550 6.700 ;
    END
  END en
  PIN sl1
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 17.250 3.450 41.000 4.050 ;
        RECT 20.000 8.450 41.000 9.050 ;
        RECT 40.400 3.450 41.000 9.050 ;
        RECT 26.450 8.400 41.000 9.050 ;
    END
  END sl1
  PIN x0
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.000 4.700 9.000 5.300 ;
    END
  END x0
  PIN x1
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.750 4.700 11.750 5.300 ;
    END
  END x1
  PIN x2
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 32.750 4.700 34.750 5.300 ;
    END
  END x2
  PIN x3
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 29.500 4.700 31.500 5.300 ;
    END
  END x3
  OBS 
      LAYER Metal1 ;
        RECT 3.700 8.400 19.350 9.000 ;
        RECT 2.650 7.200 38.600 7.800 ;
  END 
END deche4_8

MACRO deche4_4
  CLASS  CORE ;
  FOREIGN deche4_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 37.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 2.200 0.000 2.800 2.700 ;
        RECT 0.000 0.000 37.500 2.500 ;
        RECT 34.700 0.000 35.300 2.700 ;
    END
  END vss!
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 6.650 13.550 7.250 16.250 ;
        RECT 0.000 13.750 37.500 16.250 ;
        RECT 30.250 13.550 30.850 16.250 ;
    END
  END vdd!
  PIN sl0
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 18.150 8.450 20.500 9.050 ;
    END
  END sl0
  PIN en
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.050 5.950 5.850 6.550 ;
        RECT 31.650 6.100 34.650 6.700 ;
        RECT 5.250 7.200 32.250 7.800 ;
        RECT 31.650 6.100 32.250 7.800 ;
        RECT 5.250 5.950 5.850 7.800 ;
    END
  END en
  PIN sl1
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 18.150 4.700 33.350 5.300 ;
    END
  END sl1
  PIN x0
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 8.450 2.250 9.050 ;
    END
  END x0
  PIN x1
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.250 8.450 9.250 9.050 ;
    END
  END x1
  PIN x2
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 35.250 8.450 37.250 9.050 ;
    END
  END x2
  PIN x3
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 28.250 8.450 30.250 9.050 ;
    END
  END x3
  OBS 
      LAYER Metal1 ;
        RECT 1.750 7.200 4.550 7.800 ;
        RECT 9.750 8.350 10.350 9.050 ;
        RECT 9.750 8.450 16.200 9.050 ;
        RECT 4.150 4.700 17.500 5.300 ;
        RECT 27.150 8.350 27.750 9.050 ;
        RECT 21.300 8.450 27.750 9.050 ;
        RECT 6.400 5.950 31.100 6.550 ;
        RECT 32.950 7.200 35.750 7.800 ;
  END 
END deche4_4

MACRO deche4_2
  CLASS  CORE ;
  FOREIGN deche4_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 27.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 27.500 2.500 ;
    END
  END vss!
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 2.150 13.550 2.750 16.250 ;
        RECT 0.000 13.750 27.500 16.250 ;
        RECT 24.750 13.550 25.350 16.250 ;
        RECT 21.750 13.550 22.350 16.250 ;
        RECT 5.150 13.550 5.750 16.250 ;
    END
  END vdd!
  PIN sl0
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 13.850 8.350 15.550 9.150 ;
    END
  END sl0
  PIN en
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.100 3.450 20.450 4.050 ;
    END
  END en
  PIN sl1
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 13.100 5.950 20.300 6.550 ;
        RECT 19.700 5.950 20.300 7.650 ;
    END
  END sl1
  PIN x0
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.300 5.950 4.300 6.550 ;
    END
  END x0
  PIN x1
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 8.450 2.250 9.050 ;
    END
  END x1
  PIN x2
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 23.250 5.950 25.250 6.550 ;
    END
  END x2
  PIN x3
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 25.250 8.450 27.250 9.050 ;
    END
  END x3
  OBS 
      LAYER Metal1 ;
        RECT 4.750 7.800 5.350 8.750 ;
        RECT 4.750 8.150 10.850 8.750 ;
        RECT 8.000 5.950 12.400 6.550 ;
        RECT 8.000 5.950 8.600 7.650 ;
        RECT 9.150 7.050 12.400 7.650 ;
        RECT 11.800 7.200 18.400 7.800 ;
        RECT 22.200 7.800 22.800 8.900 ;
        RECT 16.650 8.300 22.800 8.900 ;
  END 
END deche4_2

MACRO deche4_1
  CLASS  CORE ;
  FOREIGN deche4_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 25.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 25.000 2.500 ;
    END
  END vss!
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 25.000 16.250 ;
    END
  END vdd!
  PIN sl0
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 12.100 8.450 14.250 9.050 ;
    END
  END sl0
  PIN en
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.600 6.850 5.300 7.800 ;
        RECT 4.600 7.200 20.600 7.800 ;
        RECT 20.000 6.750 20.600 7.800 ;
    END
  END en
  PIN sl1
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 11.800 4.700 16.550 5.300 ;
        RECT 15.950 5.950 19.300 6.550 ;
        RECT 15.950 4.700 16.550 6.550 ;
    END
  END sl1
  PIN x0
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.000 5.950 3.000 6.550 ;
    END
  END x0
  PIN x1
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 8.450 2.250 9.050 ;
    END
  END x1
  PIN x2
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 22.000 5.950 24.000 6.550 ;
    END
  END x2
  PIN x3
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 22.750 8.450 24.750 9.050 ;
    END
  END x3
  OBS 
      LAYER Metal1 ;
        RECT 3.450 8.450 9.550 9.050 ;
        RECT 6.550 4.800 11.100 5.400 ;
        RECT 6.550 4.800 7.150 6.550 ;
        RECT 5.750 5.950 7.150 6.550 ;
        RECT 7.850 6.000 14.500 6.600 ;
        RECT 15.450 8.450 21.550 9.050 ;
  END 
END deche4_1

MACRO corefill_6
  CLASS  CORE ;
  FOREIGN corefill_6 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 7.500 2.500 ;
    END
  END vss!
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 7.500 16.250 ;
    END
  END vdd!
END corefill_6

MACRO corefill_5
  CLASS  CORE ;
  FOREIGN corefill_5 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 6.250 2.500 ;
    END
  END vss!
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 6.250 16.250 ;
    END
  END vdd!
END corefill_5

MACRO corefill_4
  CLASS  CORE ;
  FOREIGN corefill_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 5.000 2.500 ;
    END
  END vss!
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 5.000 16.250 ;
    END
  END vdd!
END corefill_4

MACRO corefill_3
  CLASS  CORE ;
  FOREIGN corefill_3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 3.750 2.500 ;
    END
  END vss!
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 3.750 16.250 ;
    END
  END vdd!
END corefill_3

MACRO corefill_2
  CLASS  CORE ;
  FOREIGN corefill_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 2.500 2.500 ;
    END
  END vss!
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 2.500 16.250 ;
    END
  END vdd!
END corefill_2

MACRO corefill_1
  CLASS  CORE ;
  FOREIGN corefill_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 1.250 2.500 ;
    END
  END vss!
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 1.250 16.250 ;
    END
  END vdd!
END corefill_1

MACRO bushold
  CLASS  CORE ;
  FOREIGN bushold 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 2.050 0.000 2.650 2.650 ;
        RECT 0.000 0.000 6.250 2.500 ;
    END
  END vss!
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 2.150 13.450 2.750 16.250 ;
        RECT 0.000 13.750 6.250 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION INOUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.750 8.450 5.250 9.050 ;
    END
  END x
END bushold

MACRO buf_8
  CLASS  CORE ;
  FOREIGN buf_8 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.850 8.450 3.100 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 10.000 2.500 ;
    END
  END vss!
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 10.000 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.500 8.450 9.600 9.050 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 2.150 7.200 8.450 7.800 ;
  END 
END buf_8

MACRO buf_7
  CLASS  CORE ;
  FOREIGN buf_7 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.900 5.850 4.050 6.550 ;
        RECT 0.850 5.950 4.050 6.550 ;
        RECT 3.350 5.750 4.050 6.550 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 1.000 0.000 1.600 2.650 ;
        RECT 0.000 0.000 8.750 2.500 ;
    END
  END vss!
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 4.150 13.600 4.750 16.250 ;
        RECT 0.000 13.750 8.750 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.800 5.950 7.900 6.550 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 2.650 4.650 5.350 5.250 ;
  END 
END buf_7

MACRO buf_6
  CLASS  CORE ;
  FOREIGN buf_6 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.550 7.200 4.150 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 8.750 2.500 ;
    END
  END vss!
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 8.750 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.700 7.200 7.900 7.800 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 1.350 5.950 5.300 6.550 ;
  END 
END buf_6

MACRO buf_5
  CLASS  CORE ;
  FOREIGN buf_5 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.850 8.450 2.850 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 7.500 2.500 ;
    END
  END vss!
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 7.500 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.300 8.450 6.600 9.050 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 0.700 7.200 3.750 7.800 ;
  END 
END buf_5

MACRO buf_4
  CLASS  CORE ;
  FOREIGN buf_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.750 8.450 2.750 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 6.250 2.500 ;
    END
  END vss!
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 6.250 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.450 8.450 5.800 9.050 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 0.350 7.200 3.350 7.800 ;
  END 
END buf_4

MACRO buf_3
  CLASS  CORE ;
  FOREIGN buf_3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 8.450 2.250 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 5.000 2.500 ;
    END
  END vss!
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 5.000 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.750 8.450 4.750 9.050 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 0.350 7.200 3.450 7.800 ;
  END 
END buf_3

MACRO buf_2
  CLASS  CORE ;
  FOREIGN buf_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 8.450 2.250 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 5.000 2.500 ;
    END
  END vss!
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 5.000 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.750 8.450 4.750 9.050 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 0.450 7.050 3.450 7.650 ;
  END 
END buf_2

MACRO buf_16
  CLASS  CORE ;
  FOREIGN buf_16 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.850 7.200 4.150 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 13.750 2.500 ;
    END
  END vss!
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 13.750 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.100 5.950 9.700 7.800 ;
        RECT 5.650 7.200 13.150 7.800 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 2.300 5.950 8.600 6.550 ;
  END 
END buf_16

MACRO buf_14
  CLASS  CORE ;
  FOREIGN buf_14 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.850 8.450 4.150 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 12.500 2.500 ;
    END
  END vss!
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 12.500 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.800 8.450 10.400 9.050 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 2.450 5.950 10.950 6.550 ;
  END 
END buf_14

MACRO buf_12
  CLASS  CORE ;
  FOREIGN buf_12 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.850 7.200 4.150 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 11.250 2.500 ;
    END
  END vss!
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 11.250 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.050 8.450 9.150 9.050 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 2.150 5.950 10.350 6.550 ;
  END 
END buf_12

MACRO buf_10
  CLASS  CORE ;
  FOREIGN buf_10 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.850 8.450 4.150 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 10.000 2.500 ;
    END
  END vss!
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 10.000 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.500 8.450 9.600 9.050 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 2.150 5.950 8.450 6.550 ;
  END 
END buf_10

MACRO buf_1
  CLASS  CORE ;
  FOREIGN buf_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 8.450 2.250 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 5.000 2.500 ;
    END
  END vss!
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 5.000 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.750 8.450 4.750 9.050 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 0.450 7.050 3.450 7.650 ;
  END 
END buf_1

MACRO aoi44_6
  CLASS  CORE ;
  FOREIGN aoi44_6 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 40.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 10.300 5.950 12.450 6.750 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 40.000 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 15.100 5.950 15.700 7.800 ;
        RECT 13.000 7.200 15.700 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.950 5.950 5.600 6.550 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.850 7.200 3.750 7.800 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 21.800 5.950 24.150 6.550 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 31.500 13.500 32.200 16.250 ;
        RECT 0.000 13.750 40.000 16.250 ;
    END
  END vdd!
  PIN f
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 19.700 6.900 20.300 7.800 ;
        RECT 19.700 7.200 21.650 7.800 ;
    END
  END f
  PIN g
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 27.800 6.900 28.450 7.800 ;
        RECT 27.300 7.200 29.700 7.800 ;
    END
  END g
  PIN h
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 34.550 7.200 38.500 7.800 ;
    END
  END h
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 16.200 4.850 17.000 9.050 ;
        RECT 12.200 4.850 21.100 5.450 ;
        RECT 0.950 8.450 17.900 9.050 ;
        RECT 16.200 8.350 17.200 9.050 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 2.650 9.700 37.250 10.300 ;
  END 
END aoi44_6

MACRO aoi44_5
  CLASS  CORE ;
  FOREIGN aoi44_5 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 35.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.450 5.950 10.300 6.550 ;
        RECT 9.700 5.950 10.300 6.750 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 35.000 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 13.450 5.950 14.050 7.800 ;
        RECT 13.450 5.950 14.200 6.550 ;
        RECT 11.600 7.200 14.050 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.100 5.950 4.750 6.550 ;
        RECT 4.050 5.950 4.750 6.750 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.450 7.200 2.750 7.800 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 20.600 5.850 22.250 6.750 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 35.000 16.250 ;
    END
  END vdd!
  PIN f
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 17.150 6.900 19.150 7.800 ;
    END
  END f
  PIN g
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 25.950 6.900 26.550 7.800 ;
        RECT 25.450 7.200 27.850 7.800 ;
    END
  END g
  PIN h
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 30.800 7.200 33.250 7.800 ;
    END
  END h
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 14.700 4.850 15.300 9.050 ;
        RECT 10.700 4.850 19.300 5.450 ;
        RECT 2.700 8.450 16.450 9.050 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 1.000 9.700 32.200 10.300 ;
  END 
END aoi44_5

MACRO aoi44_4
  CLASS  CORE ;
  FOREIGN aoi44_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 31.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.450 5.950 9.050 7.950 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 31.250 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 12.250 5.950 12.900 7.800 ;
        RECT 11.600 7.200 12.900 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.200 5.950 4.850 6.550 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.850 7.200 3.550 7.800 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 18.700 5.950 20.700 6.550 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 31.250 16.250 ;
    END
  END vdd!
  PIN f
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 15.650 6.950 16.250 7.800 ;
        RECT 15.650 7.200 17.900 7.800 ;
    END
  END f
  PIN g
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 22.500 6.950 24.050 7.800 ;
    END
  END g
  PIN h
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 28.150 7.200 30.300 7.850 ;
    END
  END h
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 13.450 4.850 14.050 9.050 ;
        RECT 9.950 4.850 18.050 5.450 ;
        RECT 1.300 8.450 14.050 9.050 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 3.000 9.700 30.800 10.300 ;
  END 
END aoi44_4

MACRO aoi44_3
  CLASS  CORE ;
  FOREIGN aoi44_3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 26.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.800 5.950 8.800 6.550 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 26.250 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 10.350 5.950 11.000 7.800 ;
        RECT 9.600 7.200 11.000 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.700 5.950 4.700 6.550 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.300 8.450 2.300 9.050 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 17.100 5.950 19.100 6.550 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 16.350 13.550 17.050 16.250 ;
        RECT 0.000 13.750 26.250 16.250 ;
        RECT 23.150 13.550 23.850 16.250 ;
    END
  END vdd!
  PIN f
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 13.750 6.950 15.400 7.800 ;
    END
  END f
  PIN g
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 19.700 6.950 20.300 7.800 ;
        RECT 19.700 7.200 22.000 7.800 ;
    END
  END g
  PIN h
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 24.000 8.450 26.000 9.050 ;
    END
  END h
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 12.200 4.850 12.800 9.050 ;
        RECT 8.300 4.850 15.750 5.450 ;
        RECT 12.100 4.850 12.900 5.950 ;
        RECT 2.800 8.450 12.800 9.050 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 1.100 9.700 25.500 10.300 ;
  END 
END aoi44_3

MACRO aoi44_2
  CLASS  CORE ;
  FOREIGN aoi44_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 22.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.800 5.950 8.800 6.550 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 22.500 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.600 7.200 6.700 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.450 5.950 3.750 6.550 ;
        RECT 3.150 5.950 3.750 7.900 ;
        RECT 2.900 5.950 3.750 6.650 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.650 7.200 2.650 7.800 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 13.450 5.950 14.050 6.750 ;
        RECT 13.450 5.950 15.300 6.550 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 11.050 13.550 11.750 16.250 ;
        RECT 0.000 13.750 22.500 16.250 ;
        RECT 17.850 13.550 18.550 16.250 ;
        RECT 14.450 13.550 15.150 16.250 ;
    END
  END vdd!
  PIN f
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 10.800 6.900 11.550 7.800 ;
        RECT 10.800 7.200 12.750 7.800 ;
    END
  END f
  PIN g
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 15.950 5.950 16.550 6.750 ;
        RECT 15.950 5.950 17.900 6.550 ;
    END
  END g
  PIN h
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 19.700 8.450 21.700 9.050 ;
    END
  END h
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.350 4.700 11.700 5.300 ;
        RECT 9.700 4.700 11.700 5.450 ;
        RECT 0.850 8.450 10.300 9.050 ;
        RECT 9.700 4.700 10.300 9.050 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 2.550 9.700 20.200 10.300 ;
  END 
END aoi44_2

MACRO aoi44_1
  CLASS  CORE ;
  FOREIGN aoi44_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.450 5.950 9.050 7.950 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 15.000 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.600 7.100 11.100 7.900 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 11.650 7.200 12.250 8.550 ;
        RECT 11.650 7.200 14.550 7.800 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 12.750 8.450 14.750 9.050 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.950 5.950 6.800 6.550 ;
        RECT 6.200 5.950 6.800 8.000 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 15.000 16.250 ;
    END
  END vdd!
  PIN f
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.800 7.200 5.350 7.800 ;
        RECT 4.750 8.450 5.400 9.050 ;
        RECT 4.750 7.200 5.350 9.050 ;
    END
  END f
  PIN g
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.650 5.950 3.050 6.550 ;
        RECT 2.450 5.950 3.050 8.500 ;
    END
  END g
  PIN h
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 8.350 1.750 9.150 ;
    END
  END h
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.300 7.400 7.900 10.300 ;
        RECT 7.300 9.700 12.850 10.300 ;
        RECT 7.300 9.600 8.350 10.300 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 0.450 11.000 14.600 11.600 ;
  END 
END aoi44_1

MACRO aoi33_6
  CLASS  CORE ;
  FOREIGN aoi33_6 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 35.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 10.300 5.850 10.950 7.800 ;
        RECT 10.300 5.850 13.000 6.450 ;
        RECT 1.800 7.200 10.950 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 9.650 0.000 10.250 2.800 ;
        RECT 0.000 0.000 35.000 2.500 ;
        RECT 31.200 0.000 31.900 2.700 ;
        RECT 23.600 0.000 24.300 2.700 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.050 5.950 9.050 6.550 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 14.450 7.200 15.300 7.800 ;
        RECT 14.700 7.200 15.300 9.050 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 23.150 7.150 23.750 9.050 ;
        RECT 22.100 8.450 27.450 9.050 ;
        RECT 26.850 7.050 27.450 9.050 ;
        RECT 26.650 8.350 27.450 9.050 ;
        RECT 22.100 8.350 23.750 9.050 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 24.250 7.150 26.200 7.800 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 35.000 16.250 ;
    END
  END vdd!
  PIN f
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 24.150 5.850 25.000 6.550 ;
        RECT 17.450 5.950 30.500 6.550 ;
    END
  END f
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 20.150 3.400 27.750 4.050 ;
        RECT 5.950 3.450 27.750 4.050 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 2.750 8.450 13.550 9.050 ;
        RECT 0.900 9.700 32.300 10.300 ;
  END 
END aoi33_6

MACRO aoi33_5
  CLASS  CORE ;
  FOREIGN aoi33_5 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 31.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 12.150 6.000 12.750 7.800 ;
        RECT 0.850 7.200 12.750 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 2.050 0.000 2.650 2.750 ;
        RECT 0.000 0.000 31.250 2.500 ;
        RECT 23.450 0.000 24.050 2.700 ;
        RECT 16.400 0.000 17.100 2.700 ;
        RECT 9.250 0.000 9.850 2.700 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.050 5.750 2.650 6.550 ;
        RECT 2.050 5.950 11.650 6.550 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 13.250 7.200 16.550 7.800 ;
        RECT 15.950 7.200 16.550 9.150 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 14.300 5.950 14.900 6.600 ;
        RECT 14.300 5.950 26.800 6.550 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 20.250 7.200 23.700 7.800 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 31.250 16.250 ;
    END
  END vdd!
  PIN f
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 18.450 7.200 19.050 9.050 ;
        RECT 18.450 8.450 30.800 9.050 ;
        RECT 24.050 8.350 24.850 9.050 ;
        RECT 24.250 7.200 24.850 9.050 ;
    END
  END f
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 19.950 4.650 27.550 5.300 ;
        RECT 5.550 4.700 27.550 5.300 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 2.150 8.450 12.950 9.050 ;
        RECT 0.450 9.700 28.250 10.300 ;
        RECT 27.650 9.700 28.250 10.400 ;
  END 
END aoi33_5

MACRO aoi33_4
  CLASS  CORE ;
  FOREIGN aoi33_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 26.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.350 7.200 10.200 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 2.050 0.000 2.650 2.750 ;
        RECT 0.000 0.000 26.250 2.500 ;
        RECT 9.250 0.000 9.850 2.800 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.450 5.900 11.650 6.550 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.200 5.950 8.950 6.550 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 12.900 5.950 21.250 6.550 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 22.250 5.950 24.250 6.550 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 15.700 13.500 16.400 16.250 ;
        RECT 0.000 13.750 26.250 16.250 ;
        RECT 19.100 13.500 19.800 16.250 ;
    END
  END vdd!
  PIN f
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 14.600 7.100 15.350 7.800 ;
        RECT 14.600 7.200 25.350 7.800 ;
    END
  END f
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 19.950 4.650 20.550 5.300 ;
        RECT 5.550 4.700 20.550 5.300 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 2.150 8.450 9.600 9.050 ;
        RECT 0.450 9.700 24.850 10.300 ;
  END 
END aoi33_4

MACRO aoi33_3
  CLASS  CORE ;
  FOREIGN aoi33_3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 23.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.950 5.950 1.550 7.800 ;
        RECT 6.650 5.950 7.450 7.650 ;
        RECT 0.950 5.950 7.450 6.550 ;
        RECT 0.450 7.200 1.550 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 2.250 0.000 2.850 2.750 ;
        RECT 0.000 0.000 23.750 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.350 7.200 5.350 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.350 7.200 10.350 7.800 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 14.450 6.100 15.050 7.800 ;
        RECT 14.450 7.200 22.900 7.800 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 18.350 5.950 20.400 6.550 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 23.750 16.250 ;
    END
  END vdd!
  PIN f
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 10.850 5.950 12.250 6.550 ;
        RECT 11.650 5.950 12.250 7.850 ;
    END
  END f
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.750 3.450 20.450 4.050 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 2.100 9.700 9.550 10.300 ;
        RECT 0.450 10.900 21.450 11.500 ;
  END 
END aoi33_3

MACRO aoi33_2
  CLASS  CORE ;
  FOREIGN aoi33_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 20.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.800 7.200 2.850 7.850 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 20.000 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.450 7.200 5.500 7.850 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.050 7.200 9.100 7.800 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 15.550 7.200 17.550 7.800 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 12.950 7.200 14.950 7.800 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 14.750 13.500 15.450 16.250 ;
        RECT 0.000 13.750 20.000 16.250 ;
    END
  END vdd!
  PIN f
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.650 7.200 11.650 7.800 ;
    END
  END f
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.500 5.950 19.150 6.550 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 0.850 9.700 8.600 10.300 ;
        RECT 6.950 3.450 14.450 4.050 ;
        RECT 2.150 10.950 17.100 11.550 ;
        RECT 15.550 3.450 19.650 4.050 ;
  END 
END aoi33_2

MACRO aoi33_1
  CLASS  CORE ;
  FOREIGN aoi33_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.850 7.200 3.250 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 12.500 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.100 8.450 3.350 9.050 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.000 7.200 5.600 9.050 ;
        RECT 5.000 7.200 7.900 7.800 ;
        RECT 5.000 7.200 5.950 7.900 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.800 8.450 11.550 9.050 ;
        RECT 10.950 8.450 11.550 10.400 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.450 8.350 9.050 10.400 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 12.500 16.250 ;
    END
  END vdd!
  PIN f
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.400 8.450 7.000 10.300 ;
        RECT 5.850 9.700 7.000 10.300 ;
    END
  END f
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.850 5.950 4.450 10.250 ;
        RECT 0.450 5.950 10.700 6.550 ;
        RECT 3.850 5.950 4.700 6.650 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 2.150 10.950 9.550 11.550 ;
  END 
END aoi33_1

MACRO aoi31_6
  CLASS  CORE ;
  FOREIGN aoi31_6 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 25.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 11.150 7.200 24.550 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 13.200 0.000 13.900 2.750 ;
        RECT 0.000 0.000 25.000 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.450 7.200 10.350 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 11.550 5.900 14.000 6.550 ;
        RECT 6.400 5.950 24.100 6.550 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.750 5.950 5.600 6.550 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 10.600 13.550 11.300 16.250 ;
        RECT 0.000 13.750 25.000 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.850 3.450 17.350 4.050 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 2.150 9.700 22.850 10.300 ;
  END 
END aoi31_6

MACRO aoi31_5
  CLASS  CORE ;
  FOREIGN aoi31_5 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 22.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 12.500 7.150 15.700 7.800 ;
        RECT 0.850 7.200 15.700 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 12.900 0.000 13.600 2.700 ;
        RECT 0.000 0.000 22.500 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 16.900 7.150 20.850 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.750 5.950 19.850 6.550 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.050 5.950 5.850 6.550 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 22.500 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.950 3.450 17.100 4.050 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 2.450 9.700 20.050 10.300 ;
  END 
END aoi31_5

MACRO aoi31_4
  CLASS  CORE ;
  FOREIGN aoi31_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 18.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.800 5.950 17.800 6.550 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 4.000 0.000 4.700 2.600 ;
        RECT 0.000 0.000 18.750 2.500 ;
        RECT 11.100 0.000 11.700 2.700 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 11.750 7.200 14.050 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.600 7.200 9.150 7.850 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.850 7.200 2.900 7.800 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 18.750 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.300 4.700 15.200 5.300 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 0.600 9.700 18.200 10.300 ;
  END 
END aoi31_4

MACRO aoi31_3
  CLASS  CORE ;
  FOREIGN aoi31_3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.950 5.950 6.550 7.800 ;
        RECT 5.950 5.950 9.250 6.550 ;
        RECT 3.400 7.200 6.550 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.450 0.000 1.050 2.600 ;
        RECT 0.000 0.000 15.000 2.500 ;
        RECT 5.650 0.000 6.250 2.700 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 11.000 7.200 14.050 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.750 5.950 10.350 7.850 ;
        RECT 9.750 5.950 12.800 6.550 ;
        RECT 8.250 7.200 10.350 7.850 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 7.200 2.250 7.800 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 15.000 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.150 4.700 9.750 5.300 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 0.450 9.700 14.550 10.300 ;
  END 
END aoi31_3

MACRO aoi31_2
  CLASS  CORE ;
  FOREIGN aoi31_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.700 5.950 10.300 7.800 ;
        RECT 9.700 5.950 13.200 6.550 ;
        RECT 7.250 7.200 10.300 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 13.750 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 10.900 7.200 12.900 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.750 7.200 6.750 7.800 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.850 7.200 4.250 7.800 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 9.100 13.550 9.800 16.250 ;
        RECT 0.000 13.750 13.750 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.350 5.950 8.150 6.550 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 0.650 9.700 11.450 10.300 ;
  END 
END aoi31_2

MACRO aoi31_1
  CLASS  CORE ;
  FOREIGN aoi31_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.750 8.450 4.800 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 6.050 0.000 6.650 2.700 ;
        RECT 0.000 0.000 8.750 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.350 8.450 8.350 9.050 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.150 5.950 8.150 6.550 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.950 8.450 1.550 10.300 ;
        RECT 0.950 8.450 2.250 9.050 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 8.750 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.850 5.950 1.450 6.650 ;
        RECT 0.850 5.950 3.150 6.550 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 2.550 9.700 6.550 10.300 ;
  END 
END aoi31_1

MACRO aoi23_6
  CLASS  CORE ;
  FOREIGN aoi23_6 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 30.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.900 5.950 4.150 6.550 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 17.100 0.000 17.800 2.700 ;
        RECT 0.000 0.000 30.000 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.850 5.950 9.600 6.550 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 15.750 7.050 16.350 7.800 ;
        RECT 15.750 7.200 29.100 7.800 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 24.700 5.950 26.700 6.550 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 11.050 5.950 24.200 6.550 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 15.700 13.550 16.400 16.250 ;
        RECT 0.000 13.750 30.000 16.250 ;
        RECT 22.500 13.550 23.200 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.150 4.700 28.250 5.300 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 0.450 7.200 9.550 7.800 ;
        RECT 2.150 7.200 2.750 7.900 ;
        RECT 0.450 9.700 27.850 10.300 ;
  END 
END aoi23_6

MACRO aoi23_5
  CLASS  CORE ;
  FOREIGN aoi23_5 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 27.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.650 5.950 2.600 6.700 ;
        RECT 0.850 5.950 2.850 6.550 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 16.550 0.000 17.250 2.700 ;
        RECT 0.000 0.000 27.500 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.500 5.950 8.500 6.550 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 14.950 7.100 15.850 7.800 ;
        RECT 14.950 7.200 18.500 7.800 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 22.150 7.200 25.400 7.800 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 10.900 5.950 23.450 6.550 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 27.500 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.600 4.700 20.700 5.300 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 0.700 7.200 8.100 7.800 ;
        RECT 2.400 9.700 26.800 10.300 ;
  END 
END aoi23_5

MACRO aoi23_4
  CLASS  CORE ;
  FOREIGN aoi23_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 22.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.450 7.200 5.000 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 14.400 0.000 15.100 2.700 ;
        RECT 0.000 0.000 22.500 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.300 5.950 0.950 6.800 ;
        RECT 0.300 5.950 2.350 6.550 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 11.500 7.200 14.750 7.800 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 17.900 7.200 21.300 7.800 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.400 5.950 9.000 7.800 ;
        RECT 8.400 5.950 21.300 6.550 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 15.900 13.550 16.650 16.250 ;
        RECT 0.000 13.750 22.500 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.650 4.700 18.550 5.300 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 2.400 8.450 6.400 9.050 ;
        RECT 0.700 9.700 21.700 10.300 ;
  END 
END aoi23_4

MACRO aoi23_3
  CLASS  CORE ;
  FOREIGN aoi23_3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 18.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.400 5.950 5.500 6.550 ;
        RECT 4.850 5.950 5.500 6.700 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 18.750 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.850 5.950 2.850 6.550 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 11.050 7.150 12.500 7.800 ;
        RECT 11.050 7.200 17.800 7.800 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 15.300 5.950 15.900 6.700 ;
        RECT 14.150 5.950 16.150 6.550 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.200 5.950 13.650 6.550 ;
        RECT 12.900 5.950 13.650 6.600 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 18.750 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.050 4.700 17.950 5.300 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 2.400 8.450 6.400 9.050 ;
        RECT 0.700 9.700 18.300 10.300 ;
  END 
END aoi23_3

MACRO aoi23_2
  CLASS  CORE ;
  FOREIGN aoi23_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.450 5.950 2.450 6.550 ;
        RECT 1.650 5.950 2.450 6.700 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 15.000 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.450 5.950 5.350 6.700 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 12.750 7.200 13.500 7.850 ;
        RECT 12.100 7.200 14.600 7.800 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.350 7.200 10.400 7.800 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.200 5.950 12.700 6.550 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 7.200 13.500 7.900 16.250 ;
        RECT 0.000 13.750 15.000 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.350 4.700 11.650 5.300 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 0.350 7.200 4.450 7.800 ;
        RECT 2.150 9.700 12.850 10.300 ;
  END 
END aoi23_2

MACRO aoi23_1
  CLASS  CORE ;
  FOREIGN aoi23_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.550 8.450 3.600 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 11.250 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.050 7.200 4.050 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.400 7.200 10.450 7.800 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.700 7.200 7.850 7.800 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.650 8.450 6.650 9.050 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 11.250 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.450 4.700 10.000 5.300 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 0.450 8.500 1.050 10.300 ;
        RECT 0.450 9.700 2.750 10.300 ;
        RECT 0.450 10.950 9.100 11.550 ;
  END 
END aoi23_1

MACRO aoi22_6
  CLASS  CORE ;
  FOREIGN aoi22_6 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 23.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 13.350 5.950 16.550 6.550 ;
        RECT 15.950 5.900 21.350 6.500 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 6.300 0.000 7.000 2.700 ;
        RECT 0.000 0.000 23.750 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 12.250 5.950 12.850 7.800 ;
        RECT 12.250 7.200 22.900 7.800 ;
        RECT 17.300 7.000 21.250 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.900 5.950 7.400 6.550 ;
        RECT 3.600 5.950 7.400 6.650 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 10.150 7.000 10.750 7.800 ;
        RECT 7.900 7.200 10.750 7.800 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 15.800 13.550 16.500 16.250 ;
        RECT 0.000 13.750 23.750 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.350 3.450 20.000 4.050 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 2.250 7.200 6.300 7.800 ;
        RECT 0.550 9.700 21.550 10.300 ;
  END 
END aoi22_6

MACRO aoi22_5
  CLASS  CORE ;
  FOREIGN aoi22_5 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 20.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 13.100 5.950 17.400 6.550 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 4.500 0.000 5.200 2.700 ;
        RECT 0.000 0.000 20.000 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 10.500 6.000 11.100 7.800 ;
        RECT 10.500 7.200 19.150 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.400 5.950 5.400 6.550 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.100 5.950 9.150 6.550 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 20.000 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.850 3.450 18.250 4.050 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 0.400 7.200 7.850 7.800 ;
        RECT 2.150 9.700 19.550 10.300 ;
  END 
END aoi22_5

MACRO aoi22_4
  CLASS  CORE ;
  FOREIGN aoi22_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 17.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.900 5.950 17.100 6.550 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 2.100 0.000 2.700 2.700 ;
        RECT 0.000 0.000 17.500 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.400 6.000 9.000 7.800 ;
        RECT 8.400 7.200 16.000 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.450 5.950 2.900 6.550 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.600 5.950 7.550 6.550 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 17.500 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.650 3.450 10.850 4.050 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 2.400 7.200 6.400 7.800 ;
        RECT 0.700 9.700 14.900 10.300 ;
  END 
END aoi22_4

MACRO aoi22_3
  CLASS  CORE ;
  FOREIGN aoi22_3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.450 5.950 14.650 6.550 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 1.850 0.000 2.450 2.700 ;
        RECT 0.000 0.000 15.000 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.800 5.800 8.400 7.800 ;
        RECT 7.800 7.200 13.550 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.250 5.950 6.850 6.600 ;
        RECT 0.450 5.950 6.900 6.550 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.850 7.200 2.900 7.800 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 15.000 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.450 3.450 10.400 4.050 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 0.450 9.700 14.550 10.300 ;
  END 
END aoi22_3

MACRO aoi22_2
  CLASS  CORE ;
  FOREIGN aoi22_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.450 6.100 9.050 9.050 ;
        RECT 8.450 6.100 10.050 6.700 ;
        RECT 8.450 6.100 9.150 7.200 ;
        RECT 6.650 8.450 9.050 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 3.100 0.000 3.700 2.700 ;
        RECT 0.000 0.000 13.750 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 10.050 8.450 12.900 9.050 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.150 8.450 6.150 9.050 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.850 8.450 3.550 9.050 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 13.750 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.000 5.950 4.600 7.350 ;
        RECT 0.600 5.950 6.550 6.550 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 2.300 9.700 13.100 10.300 ;
  END 
END aoi22_2

MACRO aoi22_1
  CLASS  CORE ;
  FOREIGN aoi22_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.250 5.950 5.850 8.400 ;
        RECT 5.250 5.950 6.550 6.550 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 8.750 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.500 8.450 8.500 9.050 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.500 7.750 4.100 9.050 ;
        RECT 2.800 8.450 4.100 9.050 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 8.450 2.300 9.050 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 8.750 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.400 5.950 3.000 7.350 ;
        RECT 2.200 5.950 4.700 6.550 ;
        RECT 4.050 5.900 4.700 6.550 ;
        RECT 2.400 5.950 3.350 6.650 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 0.700 9.700 8.100 10.300 ;
  END 
END aoi22_1

MACRO aoi222_5
  CLASS  CORE ;
  FOREIGN aoi222_5 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 42.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.550 8.450 2.550 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 42.500 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.000 4.700 7.250 5.300 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 13.300 4.700 15.300 5.300 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 23.400 4.700 24.100 5.350 ;
        RECT 23.400 4.700 25.400 5.300 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 39.300 8.450 41.300 9.050 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 42.500 16.250 ;
    END
  END vdd!
  PIN f
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 31.250 4.700 33.250 5.300 ;
    END
  END f
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.550 3.450 30.450 4.050 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 22.150 8.500 26.200 9.100 ;
  END 
END aoi222_5

MACRO aoi222_4
  CLASS  CORE ;
  FOREIGN aoi222_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 36.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.900 4.700 7.950 5.300 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 36.250 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.650 8.450 2.650 9.050 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 19.250 4.700 21.250 5.300 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 10.700 4.700 12.700 5.300 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 31.750 8.450 33.750 9.050 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 23.850 13.600 24.450 16.250 ;
        RECT 0.000 13.750 36.250 16.250 ;
    END
  END vdd!
  PIN f
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 23.250 4.700 25.250 5.300 ;
    END
  END f
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.550 3.450 27.700 4.050 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 19.100 8.500 22.800 9.100 ;
  END 
END aoi222_4

MACRO aoi222_3
  CLASS  CORE ;
  FOREIGN aoi222_3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 31.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.750 4.700 7.750 5.300 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 31.250 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.550 8.450 2.550 9.050 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 15.800 4.700 17.800 5.300 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.450 4.700 11.450 5.300 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 25.500 4.700 27.500 5.300 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 23.850 13.600 24.450 16.250 ;
        RECT 0.000 13.750 31.250 16.250 ;
    END
  END vdd!
  PIN f
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 19.500 4.700 21.550 5.300 ;
    END
  END f
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.050 3.450 25.050 4.050 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 15.300 8.500 19.400 9.100 ;
  END 
END aoi222_3

MACRO aoi222_2
  CLASS  CORE ;
  FOREIGN aoi222_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 25.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.550 8.450 2.550 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 25.000 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.750 4.700 7.750 5.300 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 13.300 4.700 15.300 5.300 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 10.200 4.700 12.200 5.300 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 22.500 4.700 24.500 5.300 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 20.450 13.600 21.050 16.250 ;
        RECT 0.000 13.750 25.000 16.250 ;
    END
  END vdd!
  PIN f
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 17.000 4.700 19.000 5.300 ;
    END
  END f
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.550 3.450 20.350 4.050 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 10.200 8.500 14.300 9.100 ;
  END 
END aoi222_2

MACRO aoi222_1
  CLASS  CORE ;
  FOREIGN aoi222_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 20.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.400 8.450 5.400 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 20.000 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.550 8.450 2.550 9.050 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.450 4.700 8.450 5.300 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.050 4.700 11.050 5.300 ;
        RECT 10.300 4.700 11.050 5.350 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 17.500 4.700 19.500 5.300 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 15.400 13.600 16.000 16.250 ;
        RECT 0.000 13.750 20.000 16.250 ;
    END
  END vdd!
  PIN f
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 13.250 4.700 15.250 5.300 ;
    END
  END f
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.000 3.450 15.100 4.050 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 8.850 8.500 14.250 9.100 ;
  END 
END aoi222_1

MACRO aoi221_5
  CLASS  CORE ;
  FOREIGN aoi221_5 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 38.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.150 4.700 26.550 5.300 ;
        RECT 25.950 5.900 35.300 6.500 ;
        RECT 34.650 4.700 35.300 6.500 ;
        RECT 25.950 4.700 26.550 6.500 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 38.750 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 36.250 5.950 38.250 6.550 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.500 8.450 4.700 9.050 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 8.400 2.000 9.100 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 27.750 4.700 29.750 5.300 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 1.000 13.450 1.600 16.250 ;
        RECT 0.000 13.750 38.750 16.250 ;
        RECT 17.450 13.550 18.150 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.650 3.450 30.000 4.050 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 15.800 6.000 19.800 6.600 ;
  END 
END aoi221_5

MACRO aoi221_4
  CLASS  CORE ;
  FOREIGN aoi221_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 36.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.150 5.950 6.150 6.550 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 36.250 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 33.750 7.150 36.000 7.850 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.500 8.450 4.500 9.050 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 8.400 2.000 9.100 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 21.250 4.600 21.900 5.300 ;
        RECT 19.950 4.700 21.900 5.300 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 1.000 13.450 1.600 16.250 ;
        RECT 0.000 13.750 36.250 16.250 ;
        RECT 17.450 13.550 18.150 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 30.850 5.950 32.850 6.550 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 12.400 8.400 16.400 9.000 ;
        RECT 3.050 3.450 26.300 4.050 ;
        RECT 29.700 8.450 33.700 9.050 ;
  END 
END aoi221_4

MACRO aoi221_3
  CLASS  CORE ;
  FOREIGN aoi221_3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 31.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.650 4.700 6.650 5.300 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 31.250 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 29.000 3.450 31.000 4.050 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.550 4.700 3.550 5.300 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.400 7.200 2.400 7.800 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 15.000 4.700 17.000 5.300 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 1.000 13.450 1.600 16.250 ;
        RECT 0.000 13.750 31.250 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 17.500 3.000 18.450 4.050 ;
        RECT 4.700 3.450 22.000 4.050 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 10.800 7.000 15.000 7.600 ;
        RECT 9.100 5.900 16.700 6.500 ;
        RECT 16.100 5.900 16.700 7.300 ;
  END 
END aoi221_3

MACRO aoi221_2
  CLASS  CORE ;
  FOREIGN aoi221_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 27.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.000 4.700 10.300 5.300 ;
        RECT 20.950 4.650 25.900 5.300 ;
        RECT 9.700 5.900 21.550 6.500 ;
        RECT 20.950 4.650 21.550 6.500 ;
        RECT 9.700 4.700 10.300 6.500 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 27.500 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 25.250 7.200 27.250 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.850 4.700 2.850 5.300 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.300 7.200 2.300 7.800 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 14.250 4.700 16.250 5.300 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 1.050 13.450 1.650 16.250 ;
        RECT 0.000 13.750 27.500 16.250 ;
        RECT 26.450 13.450 27.050 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.700 3.450 21.000 4.050 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 10.150 8.100 14.150 8.700 ;
        RECT 8.450 7.000 17.200 7.600 ;
  END 
END aoi221_2

MACRO aoi221_1
  CLASS  CORE ;
  FOREIGN aoi221_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 20.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.750 7.200 4.750 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 20.000 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.250 4.700 8.450 5.300 ;
        RECT 7.800 4.700 8.450 5.350 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.700 4.700 11.700 5.300 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 16.450 7.200 18.450 7.800 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 7.200 2.250 7.800 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 15.400 13.600 16.000 16.250 ;
        RECT 0.000 13.750 20.000 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.850 3.450 12.800 4.050 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 5.400 7.200 14.300 7.800 ;
  END 
END aoi221_1

MACRO aoi21_6
  CLASS  CORE ;
  FOREIGN aoi21_6 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 18.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.700 5.950 16.550 6.550 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 2.400 0.000 3.000 2.700 ;
        RECT 0.000 0.000 18.750 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.100 5.950 9.100 6.550 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.000 5.900 3.600 6.550 ;
        RECT 3.000 5.950 5.800 6.550 ;
        RECT 5.200 5.900 5.800 6.550 ;
    END
  END c
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 10.850 13.550 11.550 16.250 ;
        RECT 0.000 13.750 18.750 16.250 ;
        RECT 14.250 13.550 14.950 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.700 3.450 15.000 4.050 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 2.400 9.700 16.600 10.300 ;
  END 
END aoi21_6

MACRO aoi21_5
  CLASS  CORE ;
  FOREIGN aoi21_5 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 17.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 12.150 7.200 15.550 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 11.900 0.000 12.500 2.700 ;
        RECT 0.000 0.000 17.500 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.850 7.200 9.150 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.900 7.200 3.500 7.850 ;
        RECT 5.300 7.200 5.950 7.850 ;
        RECT 2.900 7.200 5.950 7.800 ;
    END
  END c
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 17.500 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.800 4.700 15.100 5.300 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 2.500 9.700 16.700 10.300 ;
  END 
END aoi21_5

MACRO aoi21_4
  CLASS  CORE ;
  FOREIGN aoi21_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.650 7.200 11.650 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 15.000 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.500 7.200 8.600 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.150 7.200 2.750 8.000 ;
        RECT 2.150 7.200 4.150 7.800 ;
    END
  END c
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 15.000 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.850 4.700 5.750 5.300 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 0.450 8.600 4.450 9.200 ;
        RECT 2.150 9.700 12.950 10.300 ;
  END 
END aoi21_4

MACRO aoi21_3
  CLASS  CORE ;
  FOREIGN aoi21_3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.450 7.200 10.700 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 12.500 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.200 7.200 7.300 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.450 7.200 4.450 7.800 ;
    END
  END c
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 12.500 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.900 4.700 8.150 5.300 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 0.850 9.700 11.650 10.300 ;
  END 
END aoi21_3

MACRO aoi21_2
  CLASS  CORE ;
  FOREIGN aoi21_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.150 7.200 9.200 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 10.000 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.650 7.150 6.550 7.850 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.050 7.200 4.050 7.800 ;
    END
  END c
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 5.550 13.550 6.150 16.250 ;
        RECT 0.000 13.750 10.000 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.100 4.700 7.900 5.300 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 0.450 9.700 7.850 10.300 ;
  END 
END aoi21_2

MACRO aoi21_1
  CLASS  CORE ;
  FOREIGN aoi21_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.350 8.450 6.350 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 7.500 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.400 5.950 5.400 6.550 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.400 8.450 3.400 9.050 ;
    END
  END c
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 7.500 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.850 4.700 6.650 5.300 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 2.600 9.700 6.600 10.300 ;
  END 
END aoi21_1

MACRO aoi211_5
  CLASS  CORE ;
  FOREIGN aoi211_5 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 26.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.200 4.700 2.800 6.550 ;
        RECT 2.200 4.700 10.700 5.300 ;
        RECT 0.800 5.950 2.800 6.550 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 18.000 0.000 18.700 2.700 ;
        RECT 0.000 0.000 26.250 2.500 ;
        RECT 21.400 0.000 22.100 2.700 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.600 5.950 10.350 6.550 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 15.100 4.700 25.800 5.300 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 17.200 5.950 20.300 6.550 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 26.250 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.400 3.450 23.750 4.050 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 16.900 7.150 23.600 7.750 ;
        RECT 0.700 8.450 25.300 9.050 ;
  END 
END aoi211_5

MACRO aoi211_4
  CLASS  CORE ;
  FOREIGN aoi211_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 21.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.450 5.950 9.950 6.550 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 15.200 0.000 15.900 2.800 ;
        RECT 0.000 0.000 21.250 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.200 4.700 2.800 6.550 ;
        RECT 10.950 4.700 11.650 5.450 ;
        RECT 2.200 4.700 11.650 5.300 ;
        RECT 6.200 4.700 7.100 5.550 ;
        RECT 0.800 5.950 2.800 6.550 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 12.500 5.950 14.500 6.550 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 18.750 5.950 20.750 6.550 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 10.650 13.550 11.350 16.250 ;
        RECT 0.000 13.750 21.250 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.850 3.450 17.550 4.050 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 2.200 8.450 18.200 9.050 ;
        RECT 16.950 6.250 17.550 7.750 ;
        RECT 15.000 7.150 20.800 7.750 ;
  END 
END aoi211_4

MACRO aoi211_3
  CLASS  CORE ;
  FOREIGN aoi211_3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 21.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.850 5.950 7.850 6.550 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 21.250 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.600 5.950 2.600 6.550 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 11.500 5.950 13.500 6.550 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 19.000 5.950 21.000 6.550 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 3.850 13.550 4.550 16.250 ;
        RECT 0.000 13.750 21.250 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.450 5.950 4.050 7.800 ;
        RECT 3.450 7.200 20.800 7.800 ;
        RECT 17.850 5.850 18.450 7.800 ;
        RECT 14.150 5.850 15.050 7.800 ;
        RECT 8.850 5.900 9.600 7.800 ;
        RECT 3.450 5.950 4.250 6.550 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 2.200 8.450 18.200 9.050 ;
  END 
END aoi211_3

MACRO aoi211_2
  CLASS  CORE ;
  FOREIGN aoi211_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 17.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.750 7.200 8.750 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 17.500 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.100 7.200 4.100 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.650 7.200 12.850 7.800 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 14.600 7.200 16.600 7.800 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 2.350 13.550 3.050 16.250 ;
        RECT 0.000 13.750 17.500 16.250 ;
        RECT 9.150 13.550 9.850 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.700 7.200 5.850 7.800 ;
        RECT 5.250 8.450 14.100 9.050 ;
        RECT 13.500 8.100 14.100 9.050 ;
        RECT 5.250 7.200 5.850 9.050 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 0.700 9.700 16.700 10.300 ;
  END 
END aoi211_2

MACRO aoi211_1
  CLASS  CORE ;
  FOREIGN aoi211_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.500 7.200 7.500 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 13.750 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.600 7.200 2.600 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 10.900 7.200 12.900 7.800 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.250 7.200 10.250 7.800 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 13.750 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.450 7.200 4.600 7.800 ;
        RECT 4.000 8.450 10.700 9.050 ;
        RECT 4.000 7.200 4.600 9.050 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 0.450 9.700 13.300 10.300 ;
  END 
END aoi211_1

MACRO aoai211_5
  CLASS  CORE ;
  FOREIGN aoai211_5 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 21.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 16.100 5.900 16.700 6.550 ;
        RECT 11.200 5.950 16.700 6.550 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 5.650 0.000 6.250 2.800 ;
        RECT 0.000 0.000 21.250 2.500 ;
        RECT 13.850 0.000 14.450 2.800 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.500 7.200 19.900 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.850 7.200 5.850 7.800 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.650 7.200 2.650 7.800 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 21.250 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.450 9.700 7.850 10.300 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 0.450 4.700 17.050 5.300 ;
        RECT 8.950 9.700 19.750 10.300 ;
  END 
END aoai211_5

MACRO aoai211_4
  CLASS  CORE ;
  FOREIGN aoai211_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 18.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.100 5.950 8.700 7.800 ;
        RECT 8.100 7.200 18.150 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 5.650 0.000 6.250 2.800 ;
        RECT 0.000 0.000 18.750 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 14.150 5.900 15.000 6.550 ;
        RECT 9.500 5.950 15.000 6.550 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.950 5.950 6.950 6.550 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.650 7.200 2.650 7.800 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.450 13.450 1.050 16.250 ;
        RECT 0.000 13.750 18.750 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.150 9.700 7.450 10.300 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 0.450 4.700 13.150 5.300 ;
        RECT 8.550 9.700 15.950 10.300 ;
  END 
END aoai211_4

MACRO aoai211_3
  CLASS  CORE ;
  FOREIGN aoai211_3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 16.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 13.850 8.450 15.050 9.100 ;
        RECT 13.850 8.450 15.800 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 5.650 0.000 6.250 2.800 ;
        RECT 0.000 0.000 16.250 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.100 7.200 14.350 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.800 7.200 6.800 7.800 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.500 7.200 2.500 7.800 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 10.050 13.500 10.750 16.250 ;
        RECT 0.000 13.750 16.250 16.250 ;
        RECT 13.450 13.500 14.150 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.150 9.700 7.300 10.300 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 0.450 3.450 11.950 4.050 ;
        RECT 8.400 9.700 15.800 10.300 ;
  END 
END aoai211_3

MACRO aoai211_2
  CLASS  CORE ;
  FOREIGN aoai211_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.150 8.450 10.150 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 5.450 0.000 6.050 2.800 ;
        RECT 0.000 0.000 12.500 2.500 ;
        RECT 10.700 0.000 11.300 2.800 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.400 5.950 11.900 6.550 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.500 5.950 4.100 7.800 ;
        RECT 3.500 7.200 11.900 7.800 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.500 7.200 2.550 7.800 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 6.100 13.500 6.800 16.250 ;
        RECT 0.000 13.750 12.500 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.400 9.700 3.400 10.300 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 4.450 9.700 8.600 10.300 ;
        RECT 0.350 3.450 8.750 4.050 ;
  END 
END aoai211_2

MACRO aoai211_1
  CLASS  CORE ;
  FOREIGN aoai211_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.450 5.950 8.450 6.550 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 3.850 0.000 4.450 2.800 ;
        RECT 0.000 0.000 10.000 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.850 7.200 6.900 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.150 8.450 5.400 9.050 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.500 7.200 2.500 7.800 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 10.000 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.350 9.700 3.650 10.300 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 2.150 4.700 7.150 5.300 ;
        RECT 4.750 9.700 8.900 10.300 ;
  END 
END aoai211_1

MACRO ao44_6
  CLASS  CORE ;
  FOREIGN ao44_6 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 30.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 21.700 7.600 22.400 9.300 ;
        RECT 21.700 8.700 29.500 9.300 ;
        RECT 21.700 8.450 22.800 9.300 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 30.000 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 28.450 7.200 29.050 8.200 ;
        RECT 25.000 7.600 29.050 8.200 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 20.650 5.950 25.350 6.550 ;
        RECT 24.750 6.500 27.800 7.100 ;
        RECT 27.200 5.850 27.800 7.100 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 18.650 4.700 19.250 6.400 ;
        RECT 25.950 4.700 26.550 6.000 ;
        RECT 18.650 4.700 26.550 5.300 ;
        RECT 18.650 4.700 19.600 5.400 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.350 8.500 0.950 9.300 ;
        RECT 0.350 8.700 8.200 9.300 ;
        RECT 7.500 7.600 8.200 9.300 ;
        RECT 7.200 8.450 8.200 9.300 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 30.000 16.250 ;
    END
  END vdd!
  PIN f
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.950 7.200 1.550 8.000 ;
        RECT 0.950 7.400 3.500 8.000 ;
    END
  END f
  PIN g
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.050 6.300 5.300 6.900 ;
        RECT 8.450 5.950 9.050 7.100 ;
        RECT 4.700 5.950 9.050 6.550 ;
    END
  END g
  PIN h
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.100 4.700 3.700 5.800 ;
        RECT 10.300 4.700 11.150 6.000 ;
        RECT 3.100 4.700 11.150 5.300 ;
    END
  END h
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 14.350 6.750 14.950 10.300 ;
        RECT 12.400 9.700 16.650 10.300 ;
        RECT 12.400 9.600 14.950 10.300 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 10.950 6.750 12.500 7.350 ;
        RECT 10.950 6.750 11.550 10.400 ;
        RECT 2.450 9.800 11.550 10.400 ;
        RECT 17.150 6.750 17.750 10.400 ;
        RECT 17.150 9.800 26.850 10.400 ;
  END 
END ao44_6

MACRO ao44_5
  CLASS  CORE ;
  FOREIGN ao44_5 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 25.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 16.700 4.700 17.300 7.150 ;
        RECT 16.700 4.700 18.200 5.300 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 25.000 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 18.950 5.950 19.600 8.000 ;
        RECT 18.950 5.950 23.450 6.550 ;
        RECT 22.800 5.800 23.450 6.550 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 20.200 7.200 20.850 9.050 ;
        RECT 20.200 7.200 24.650 7.800 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 21.750 8.450 24.400 9.050 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.450 4.650 1.250 5.300 ;
        RECT 8.050 4.700 8.650 7.150 ;
        RECT 7.900 4.700 8.650 5.400 ;
        RECT 0.450 4.700 8.650 5.300 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 2.100 13.450 2.800 16.250 ;
        RECT 0.000 13.750 25.000 16.250 ;
        RECT 22.100 13.450 22.800 16.250 ;
        RECT 12.300 13.450 13.000 16.250 ;
    END
  END vdd!
  PIN f
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.900 5.950 6.600 6.550 ;
        RECT 6.000 5.950 6.600 8.400 ;
    END
  END f
  PIN g
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.350 7.200 4.600 7.800 ;
    END
  END g
  PIN h
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.350 8.450 2.950 9.050 ;
    END
  END h
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 12.350 5.950 12.950 10.300 ;
        RECT 10.400 9.700 14.650 10.300 ;
        RECT 12.350 9.600 13.350 10.300 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 9.900 5.950 10.500 8.250 ;
        RECT 8.950 7.650 10.500 8.250 ;
        RECT 8.950 7.650 9.550 10.300 ;
        RECT 0.450 9.700 9.550 10.300 ;
        RECT 13.700 5.950 16.200 6.550 ;
        RECT 15.600 5.950 16.200 10.300 ;
        RECT 15.600 9.700 24.450 10.300 ;
  END 
END ao44_5

MACRO ao44_4
  CLASS  CORE ;
  FOREIGN ao44_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 22.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 20.900 4.650 21.500 5.300 ;
        RECT 17.800 4.700 21.500 5.300 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 22.500 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 18.650 7.000 19.700 7.800 ;
        RECT 18.650 7.200 21.950 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 16.450 7.700 17.100 9.050 ;
        RECT 16.450 8.450 22.050 9.050 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 13.550 5.950 15.000 6.600 ;
        RECT 13.550 5.950 16.800 6.550 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.400 5.950 2.450 6.550 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 22.500 16.250 ;
    END
  END vdd!
  PIN f
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.500 7.200 2.800 7.800 ;
        RECT 2.200 7.100 4.850 7.700 ;
    END
  END f
  PIN g
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.700 8.200 5.500 9.050 ;
        RECT 0.400 8.450 5.500 9.050 ;
    END
  END g
  PIN h
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.450 4.650 1.050 5.300 ;
        RECT 7.350 4.700 7.950 7.050 ;
        RECT 0.450 4.700 7.950 5.300 ;
    END
  END h
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.700 9.700 13.950 10.300 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 3.350 5.950 6.850 6.550 ;
        RECT 6.250 5.950 6.850 8.250 ;
        RECT 6.250 7.650 9.600 8.250 ;
        RECT 8.350 7.650 8.950 10.300 ;
        RECT 2.950 9.700 8.950 10.300 ;
        RECT 10.350 7.650 15.700 8.250 ;
        RECT 15.100 7.650 15.700 10.300 ;
        RECT 15.100 9.700 20.400 10.300 ;
  END 
END ao44_4

MACRO ao44_3
  CLASS  CORE ;
  FOREIGN ao44_3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 18.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 12.000 4.700 12.600 8.000 ;
        RECT 12.000 4.700 18.050 5.300 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 16.050 0.000 16.750 2.700 ;
        RECT 0.000 0.000 18.750 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 13.150 8.450 13.800 9.100 ;
        RECT 13.150 8.450 16.600 9.050 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 13.550 7.200 15.550 7.800 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 16.400 5.950 18.400 6.550 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.600 4.650 1.250 5.300 ;
        RECT 0.600 4.700 4.150 5.300 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 10.600 13.400 11.300 16.250 ;
        RECT 0.000 13.750 18.750 16.250 ;
        RECT 14.050 13.450 14.650 16.250 ;
    END
  END vdd!
  PIN f
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.600 7.200 4.050 7.800 ;
    END
  END f
  PIN g
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.450 8.450 5.650 9.050 ;
    END
  END g
  PIN h
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.400 5.950 6.700 6.550 ;
    END
  END h
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 10.400 5.000 11.000 7.800 ;
        RECT 8.950 7.200 11.000 7.800 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 7.850 6.800 8.450 10.300 ;
        RECT 2.150 9.700 8.450 10.300 ;
        RECT 12.350 9.700 16.350 10.300 ;
  END 
END ao44_3

MACRO ao44_2
  CLASS  CORE ;
  FOREIGN ao44_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 18.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 11.550 4.700 12.150 8.000 ;
        RECT 11.550 4.700 18.350 5.300 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 18.750 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 12.950 8.450 14.050 9.100 ;
        RECT 12.950 8.450 17.650 9.050 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 13.600 7.200 17.950 7.800 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 14.950 5.950 18.400 6.550 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.850 4.700 4.550 5.300 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 18.750 16.250 ;
    END
  END vdd!
  PIN f
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.600 7.200 4.050 7.800 ;
    END
  END f
  PIN g
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.450 8.450 5.650 9.050 ;
    END
  END g
  PIN h
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.300 5.950 6.450 6.650 ;
        RECT 0.500 5.950 6.550 6.550 ;
        RECT 5.850 5.950 6.450 7.800 ;
    END
  END h
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 10.400 5.200 11.000 7.800 ;
        RECT 8.950 7.200 11.000 7.800 ;
    END
  END x
END ao44_2

MACRO ao44_1
  CLASS  CORE ;
  FOREIGN ao44_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.600 5.950 10.200 7.700 ;
        RECT 9.600 5.950 11.000 6.550 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.800 0.000 1.400 2.800 ;
        RECT 0.000 0.000 15.000 2.500 ;
        RECT 14.050 0.000 14.650 2.800 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 10.600 8.450 14.200 9.050 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 11.600 7.200 13.600 7.800 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 12.600 4.700 14.600 5.300 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.450 5.950 5.300 6.550 ;
        RECT 4.700 5.950 5.300 7.800 ;
        RECT 4.400 7.200 5.000 9.050 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 15.000 16.250 ;
    END
  END vdd!
  PIN f
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.400 8.450 3.300 9.050 ;
    END
  END f
  PIN g
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.550 7.200 2.550 7.800 ;
    END
  END g
  PIN h
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.350 4.700 4.150 5.300 ;
    END
  END h
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.600 7.200 8.600 7.800 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 5.700 8.450 6.300 10.300 ;
        RECT 3.600 9.700 6.300 10.300 ;
        RECT 8.300 8.450 8.900 10.300 ;
        RECT 8.300 9.700 11.000 10.300 ;
  END 
END ao44_1

MACRO ao33_6
  CLASS  CORE ;
  FOREIGN ao33_6 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 26.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 18.300 7.200 18.900 9.050 ;
        RECT 18.300 8.450 25.900 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 26.250 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 22.700 7.200 25.000 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 16.850 5.950 23.700 6.550 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.350 7.200 6.950 9.050 ;
        RECT 0.350 8.450 6.950 9.050 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.400 7.200 3.350 7.800 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 5.500 13.450 6.200 16.250 ;
        RECT 0.000 13.750 26.250 16.250 ;
        RECT 19.100 13.450 19.800 16.250 ;
    END
  END vdd!
  PIN f
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.800 5.950 9.200 6.550 ;
        RECT 8.550 5.950 9.200 6.800 ;
    END
  END f
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 12.200 6.750 12.800 10.300 ;
        RECT 10.400 9.700 14.650 10.300 ;
        RECT 12.200 6.750 12.950 7.400 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 5.850 4.700 10.500 5.300 ;
        RECT 9.900 4.700 10.500 8.450 ;
        RECT 8.950 7.850 10.500 8.450 ;
        RECT 8.950 7.850 9.550 10.300 ;
        RECT 0.450 9.700 9.550 10.300 ;
        RECT 14.550 4.700 20.350 5.300 ;
        RECT 14.550 4.700 15.150 9.000 ;
        RECT 15.150 8.400 15.750 10.300 ;
        RECT 15.150 9.700 24.850 10.300 ;
  END 
END ao33_6

MACRO ao33_5
  CLASS  CORE ;
  FOREIGN ao33_5 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 23.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 18.950 5.950 23.250 6.550 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 23.750 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 20.550 8.450 22.550 9.050 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 15.450 5.950 16.050 7.800 ;
        RECT 15.450 7.200 23.200 7.800 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.350 6.700 2.800 7.300 ;
        RECT 2.200 7.200 4.550 7.800 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.300 8.450 2.300 9.050 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 23.750 16.250 ;
    END
  END vdd!
  PIN f
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.150 4.700 9.300 5.350 ;
        RECT 8.700 4.700 9.300 5.600 ;
    END
  END f
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.650 9.700 13.650 10.300 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 9.800 7.000 10.400 9.050 ;
        RECT 2.850 8.450 10.400 9.050 ;
        RECT 2.850 8.450 3.450 9.250 ;
        RECT 11.950 4.700 18.800 5.300 ;
        RECT 11.950 4.700 12.550 9.050 ;
        RECT 11.950 8.450 20.050 9.050 ;
  END 
END ao33_5

MACRO ao33_4
  CLASS  CORE ;
  FOREIGN ao33_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 20.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.550 8.450 2.550 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 20.000 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.500 5.950 5.250 6.550 ;
        RECT 4.550 7.150 5.250 7.800 ;
        RECT 4.650 5.950 5.250 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.500 4.650 1.100 5.300 ;
        RECT 5.950 4.700 6.550 6.550 ;
        RECT 0.500 4.700 6.550 5.300 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 14.700 4.700 15.600 5.300 ;
        RECT 15.000 4.700 15.600 6.600 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 13.700 6.450 14.300 7.800 ;
        RECT 13.700 7.200 17.100 7.800 ;
        RECT 13.700 7.100 14.600 7.800 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 20.000 16.250 ;
    END
  END vdd!
  PIN f
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 17.700 5.950 19.700 6.550 ;
    END
  END f
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 10.200 8.600 10.800 10.300 ;
        RECT 9.550 9.700 10.800 10.300 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 1.700 7.200 3.800 7.800 ;
        RECT 3.200 7.200 3.800 9.050 ;
        RECT 8.400 6.350 9.000 9.050 ;
        RECT 3.200 8.450 9.000 9.050 ;
        RECT 11.500 6.100 12.100 9.050 ;
        RECT 11.500 8.450 17.600 9.050 ;
  END 
END ao33_4

MACRO ao33_3
  CLASS  CORE ;
  FOREIGN ao33_3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 16.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.400 5.950 2.400 6.550 ;
        RECT 1.650 5.950 2.400 6.650 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 16.250 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.250 7.200 4.250 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.800 5.950 6.800 6.650 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 13.850 5.950 14.700 6.650 ;
        RECT 13.850 5.950 15.850 6.550 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 12.900 8.450 14.900 9.050 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 16.250 16.250 ;
    END
  END vdd!
  PIN f
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.950 5.950 11.950 6.550 ;
        RECT 11.200 5.950 11.950 6.650 ;
    END
  END f
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.850 5.950 8.450 10.300 ;
        RECT 7.850 9.700 9.100 10.300 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 5.700 8.100 6.300 9.050 ;
        RECT 0.400 8.450 6.300 9.050 ;
        RECT 9.500 7.200 15.850 7.800 ;
        RECT 11.800 7.200 12.400 8.950 ;
  END 
END ao33_3

MACRO ao33_2
  CLASS  CORE ;
  FOREIGN ao33_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 12.100 7.200 14.600 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 15.000 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 10.650 5.950 12.700 6.550 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.450 8.450 11.650 9.050 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.400 8.450 2.450 9.050 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.150 7.200 4.150 7.800 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 15.000 16.250 ;
    END
  END vdd!
  PIN f
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.650 5.950 6.650 6.550 ;
    END
  END f
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.850 8.450 8.250 9.050 ;
    END
  END x
END ao33_2

MACRO ao33_1
  CLASS  CORE ;
  FOREIGN ao33_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.350 5.950 10.600 6.550 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 4.350 0.000 4.950 2.950 ;
        RECT 0.000 0.000 12.500 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.600 4.700 10.600 5.300 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 10.200 7.200 12.250 7.800 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.300 5.950 4.300 6.550 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.900 7.200 2.900 7.800 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 12.500 16.250 ;
    END
  END vdd!
  PIN f
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.450 3.450 2.900 4.050 ;
    END
  END f
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.150 7.200 8.150 7.800 ;
    END
  END x
END ao33_1

MACRO ao31_6
  CLASS  CORE ;
  FOREIGN ao31_6 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 22.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.100 7.200 10.100 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 22.500 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.400 7.200 6.400 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.500 7.200 3.500 7.800 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 19.300 8.450 21.300 9.050 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 10.900 13.550 11.600 16.250 ;
        RECT 0.000 13.750 22.500 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 12.600 12.200 16.700 12.800 ;
    END
  END x
END ao31_6

MACRO ao31_5
  CLASS  CORE ;
  FOREIGN ao31_5 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 20.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.750 5.850 8.450 6.550 ;
        RECT 7.750 5.950 9.750 6.550 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 20.000 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.850 7.200 5.850 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.700 8.450 2.700 9.050 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 17.750 8.450 19.750 9.050 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 7.350 13.600 7.950 16.250 ;
        RECT 0.000 13.750 20.000 16.250 ;
        RECT 15.400 13.550 16.200 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 10.300 12.200 14.400 12.800 ;
    END
  END x
END ao31_5

MACRO ao31_4
  CLASS  CORE ;
  FOREIGN ao31_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 17.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.450 7.200 3.450 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 17.500 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.200 7.200 6.200 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.700 5.700 7.350 6.550 ;
        RECT 6.700 5.950 8.700 6.550 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 14.650 7.200 16.650 7.800 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 7.450 13.500 8.150 16.250 ;
        RECT 0.000 13.750 17.500 16.250 ;
        RECT 10.900 13.500 11.600 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.200 12.200 13.300 12.800 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 2.350 12.200 6.450 12.800 ;
  END 
END ao31_4

MACRO ao31_3
  CLASS  CORE ;
  FOREIGN ao31_3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 8.450 2.250 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 13.750 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.100 5.950 3.100 6.550 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.850 7.200 5.850 7.800 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 10.400 7.200 12.400 7.800 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 13.750 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.300 6.700 9.050 7.300 ;
        RECT 8.450 8.450 9.550 9.050 ;
        RECT 8.450 6.700 9.050 9.050 ;
    END
  END x
END ao31_3

MACRO ao31_2
  CLASS  CORE ;
  FOREIGN ao31_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 8.450 2.250 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 12.500 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.100 5.950 3.100 6.550 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.200 5.950 6.200 6.550 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.100 8.450 11.100 9.050 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 5.900 13.550 6.600 16.250 ;
        RECT 0.000 13.750 12.500 16.250 ;
        RECT 9.300 13.550 10.000 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.200 5.850 7.800 8.200 ;
        RECT 7.200 7.600 8.250 8.200 ;
    END
  END x
END ao31_2

MACRO ao31_1
  CLASS  CORE ;
  FOREIGN ao31_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.400 5.950 2.400 6.550 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 4.800 0.000 5.400 2.700 ;
        RECT 0.000 0.000 10.000 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.900 8.450 2.900 9.050 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.600 7.200 4.600 7.800 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.100 7.200 7.100 7.800 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 10.000 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.600 7.200 9.600 7.800 ;
    END
  END x
END ao31_1

MACRO ao23_6
  CLASS  CORE ;
  FOREIGN ao23_6 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 23.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 20.550 7.200 22.550 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 23.750 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 17.650 7.200 19.650 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.050 7.200 7.050 7.800 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.300 8.350 1.800 9.150 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.900 4.700 10.900 5.300 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 23.750 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 12.450 8.450 16.550 9.050 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 11.350 7.200 15.800 7.800 ;
        RECT 11.350 7.200 11.950 9.100 ;
        RECT 2.300 8.500 11.950 9.100 ;
        RECT 12.250 4.700 19.950 5.300 ;
        RECT 12.250 4.700 12.850 5.500 ;
        RECT 15.950 4.700 16.550 5.500 ;
        RECT 19.300 8.500 23.400 9.100 ;
  END 
END ao23_6

MACRO ao23_5
  CLASS  CORE ;
  FOREIGN ao23_5 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 21.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 18.950 7.200 20.950 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 21.250 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 15.850 7.200 17.850 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.350 4.650 2.800 5.250 ;
        RECT 2.200 5.950 4.150 6.550 ;
        RECT 2.200 4.650 2.800 6.550 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.950 5.900 1.550 8.000 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.250 5.950 10.250 6.550 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 21.250 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 10.900 5.950 12.900 6.550 ;
        RECT 10.850 8.450 15.950 9.050 ;
        RECT 14.650 5.750 15.250 9.050 ;
        RECT 12.300 5.750 15.250 6.350 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 13.500 6.850 14.100 7.800 ;
        RECT 2.750 7.200 14.100 7.800 ;
        RECT 10.600 4.650 19.600 5.250 ;
  END 
END ao23_5

MACRO ao23_4
  CLASS  CORE ;
  FOREIGN ao23_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 16.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 13.900 7.200 15.900 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 16.250 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 11.950 5.950 13.950 6.550 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 8.450 2.250 9.050 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.400 5.750 4.550 6.350 ;
        RECT 3.950 5.750 4.550 7.900 ;
        RECT 3.450 5.750 4.550 6.550 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.400 4.600 6.550 5.200 ;
        RECT 5.950 7.200 6.900 7.800 ;
        RECT 5.950 4.600 6.550 7.800 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 14.550 13.650 15.350 16.250 ;
        RECT 0.000 13.750 16.250 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.500 7.200 10.150 9.050 ;
        RECT 9.500 8.450 11.650 9.050 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 7.450 6.100 9.100 6.700 ;
        RECT 1.800 6.850 2.400 7.800 ;
        RECT 1.800 7.200 3.350 7.800 ;
        RECT 2.750 7.200 3.350 9.150 ;
        RECT 7.450 6.100 8.050 9.150 ;
        RECT 2.750 8.550 8.050 9.150 ;
        RECT 10.650 6.050 11.450 6.700 ;
        RECT 10.650 6.050 11.300 7.800 ;
        RECT 10.650 7.200 13.300 7.800 ;
        RECT 12.700 7.200 13.300 9.050 ;
        RECT 12.700 8.450 15.900 9.050 ;
  END 
END ao23_4

MACRO ao23_3
  CLASS  CORE ;
  FOREIGN ao23_3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 12.450 8.450 14.450 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 15.000 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 10.200 7.200 12.200 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.950 7.100 1.550 9.150 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.450 6.050 4.050 8.050 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.000 5.950 7.000 6.550 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 15.000 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.200 7.200 9.600 7.800 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 0.450 5.800 2.750 6.400 ;
        RECT 2.150 5.800 2.750 9.150 ;
        RECT 2.150 8.550 6.200 9.150 ;
  END 
END ao23_3

MACRO ao23_2
  CLASS  CORE ;
  FOREIGN ao23_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 11.100 8.450 13.100 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 13.750 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.050 7.200 11.050 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.650 8.450 6.650 9.050 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.150 7.200 4.150 7.800 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.550 8.450 2.550 9.050 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 13.750 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.750 6.350 6.350 7.800 ;
        RECT 5.750 7.200 8.100 7.800 ;
    END
  END x
END ao23_2

MACRO ao23_1
  CLASS  CORE ;
  FOREIGN ao23_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 11.100 8.450 13.100 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 13.750 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.050 7.200 11.050 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.050 8.450 7.050 9.050 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.150 7.200 4.150 7.800 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.550 8.450 2.550 9.050 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 13.750 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.750 7.050 6.350 7.800 ;
        RECT 5.750 7.200 8.100 7.800 ;
    END
  END x
END ao23_1

MACRO ao22_6
  CLASS  CORE ;
  FOREIGN ao22_6 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 20.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.450 5.950 3.000 6.550 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 18.100 0.000 18.700 2.800 ;
        RECT 0.000 0.000 20.000 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.000 4.700 4.150 5.300 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 14.700 5.950 15.300 6.650 ;
        RECT 14.700 6.050 19.600 6.650 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 15.600 4.700 19.650 5.300 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 20.000 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.700 5.650 11.550 6.250 ;
        RECT 8.300 8.450 12.700 9.050 ;
        RECT 10.950 5.650 11.550 9.050 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 1.900 7.200 8.550 7.800 ;
        RECT 13.050 7.200 19.500 7.800 ;
  END 
END ao22_6

MACRO ao22_5
  CLASS  CORE ;
  FOREIGN ao22_5 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 18.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.000 8.450 3.550 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 18.750 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.050 5.950 5.800 6.550 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 15.550 4.700 18.150 5.300 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 12.950 5.950 15.500 6.550 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 18.750 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.050 9.700 11.450 10.300 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 2.750 7.200 6.750 7.800 ;
        RECT 11.650 5.950 12.250 7.800 ;
        RECT 11.650 7.200 16.550 7.800 ;
  END 
END ao22_5

MACRO ao22_4
  CLASS  CORE ;
  FOREIGN ao22_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 16.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.200 8.450 3.750 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 16.250 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.100 5.950 6.650 6.550 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 14.000 7.200 16.000 7.800 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.500 5.950 15.900 6.550 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 16.250 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.700 9.700 10.100 10.300 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 7.200 6.800 7.800 7.800 ;
        RECT 1.300 7.200 7.800 7.800 ;
        RECT 9.400 7.200 13.500 7.800 ;
  END 
END ao22_4

MACRO ao22_3
  CLASS  CORE ;
  FOREIGN ao22_3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.100 8.450 9.550 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 12.500 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.600 7.200 11.650 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.400 5.950 3.750 6.550 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.850 7.200 5.400 7.800 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 12.500 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.100 9.700 6.650 10.300 ;
    END
  END x
END ao22_3

MACRO ao22_2
  CLASS  CORE ;
  FOREIGN ao22_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.800 8.450 8.850 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 11.250 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.350 7.200 10.750 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.400 5.950 3.750 6.550 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.750 7.200 5.400 7.800 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 6.900 13.550 7.600 16.250 ;
        RECT 0.000 13.750 11.250 16.250 ;
        RECT 10.200 13.450 10.800 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.800 9.700 6.350 10.300 ;
    END
  END x
END ao22_2

MACRO ao22_1
  CLASS  CORE ;
  FOREIGN ao22_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.800 3.450 3.600 4.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 5.500 0.000 6.100 3.900 ;
        RECT 0.000 0.000 10.000 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.300 5.950 2.300 6.550 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.100 3.450 9.100 4.050 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.350 7.200 9.600 7.800 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 10.000 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.800 6.400 5.300 7.000 ;
        RECT 4.500 6.400 5.300 7.800 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 1.000 8.450 3.800 9.050 ;
        RECT 5.800 8.450 8.500 9.050 ;
  END 
END ao22_1

MACRO ao222_5
  CLASS  CORE ;
  FOREIGN ao222_5 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 26.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 23.850 7.200 25.850 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 3.050 0.000 3.650 2.750 ;
        RECT 0.000 0.000 26.250 2.500 ;
        RECT 22.600 0.000 23.200 2.750 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 21.100 7.200 23.100 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 15.250 7.200 17.250 7.800 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 18.450 7.150 20.350 7.850 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 7.200 2.250 7.800 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 2.700 13.500 3.300 16.250 ;
        RECT 0.000 13.750 26.250 16.250 ;
        RECT 23.350 13.500 24.050 16.250 ;
        RECT 19.950 13.550 20.650 16.250 ;
        RECT 16.550 12.900 17.200 16.250 ;
        RECT 12.850 13.550 13.600 16.250 ;
        RECT 6.050 13.550 6.750 16.250 ;
    END
  END vdd!
  PIN f
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.250 7.200 5.250 7.800 ;
    END
  END f
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.500 7.200 11.850 7.800 ;
    END
  END x
END ao222_5

MACRO ao222_4
  CLASS  CORE ;
  FOREIGN ao222_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 21.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 7.200 2.250 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 3.050 0.000 3.650 2.750 ;
        RECT 0.000 0.000 21.250 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.900 7.000 4.750 7.800 ;
        RECT 2.750 7.200 4.750 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 19.000 7.200 21.000 7.800 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 16.700 7.000 17.350 7.800 ;
        RECT 16.500 7.200 18.500 7.800 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 11.050 7.200 13.050 7.800 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 4.350 13.550 5.050 16.250 ;
        RECT 0.000 13.750 21.250 16.250 ;
        RECT 14.600 13.550 15.300 16.250 ;
        RECT 11.250 13.450 11.850 16.250 ;
        RECT 7.750 13.550 8.450 16.250 ;
    END
  END vdd!
  PIN f
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 14.500 7.000 15.100 7.800 ;
        RECT 13.850 7.200 15.900 7.800 ;
    END
  END f
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.950 8.450 10.300 9.050 ;
    END
  END x
END ao222_4

MACRO ao222_3
  CLASS  CORE ;
  FOREIGN ao222_3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 20.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.750 7.200 2.750 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 3.050 0.000 3.650 2.750 ;
        RECT 0.000 0.000 20.000 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.250 7.200 5.250 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 16.750 7.200 18.750 7.800 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 15.000 4.700 17.300 5.300 ;
        RECT 16.550 4.700 17.300 5.600 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 10.900 7.150 12.850 7.850 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 4.350 13.550 5.050 16.250 ;
        RECT 0.000 13.750 20.000 16.250 ;
        RECT 17.650 13.550 18.250 16.250 ;
        RECT 10.850 13.450 11.450 16.250 ;
        RECT 7.750 13.550 8.450 16.250 ;
    END
  END vdd!
  PIN f
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 13.450 7.200 15.550 7.800 ;
    END
  END f
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.100 7.200 10.150 7.800 ;
    END
  END x
END ao222_3

MACRO ao222_2
  CLASS  CORE ;
  FOREIGN ao222_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 18.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.650 7.200 2.700 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 18.750 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.250 7.200 5.300 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 16.100 7.200 18.250 7.800 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 14.650 4.700 16.800 5.300 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 10.100 7.200 12.700 7.800 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 4.350 13.550 5.050 16.250 ;
        RECT 0.000 13.750 18.750 16.250 ;
        RECT 10.850 13.450 11.450 16.250 ;
        RECT 7.750 13.550 8.450 16.250 ;
    END
  END vdd!
  PIN f
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 13.400 7.150 15.350 7.850 ;
    END
  END f
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.100 8.450 10.150 9.050 ;
    END
  END x
END ao222_2

MACRO ao222_1
  CLASS  CORE ;
  FOREIGN ao222_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 16.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.450 9.700 3.450 10.300 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 16.250 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.300 7.200 2.300 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 13.800 8.450 15.800 9.050 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 12.150 9.700 14.150 10.300 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.100 9.700 11.100 10.300 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 3.900 13.550 4.600 16.250 ;
        RECT 0.000 13.750 16.250 16.250 ;
        RECT 8.300 13.450 8.900 16.250 ;
        RECT 6.500 13.550 7.200 16.250 ;
    END
  END vdd!
  PIN f
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.950 7.200 11.950 7.800 ;
    END
  END f
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.850 8.450 8.900 9.050 ;
    END
  END x
END ao222_1

MACRO ao221_5
  CLASS  CORE ;
  FOREIGN ao221_5 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 23.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 21.400 7.200 23.400 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 23.750 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 18.900 7.200 20.900 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 13.250 7.200 15.250 7.800 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 16.400 7.200 18.400 7.800 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.400 7.200 2.400 7.800 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 3.850 13.550 4.550 16.250 ;
        RECT 0.000 13.750 23.750 16.250 ;
        RECT 20.650 13.500 21.350 16.250 ;
        RECT 17.250 13.550 17.950 16.250 ;
        RECT 13.850 12.900 14.500 16.250 ;
        RECT 10.700 13.550 11.400 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.250 7.200 9.650 7.800 ;
    END
  END x
END ao221_5

MACRO ao221_4
  CLASS  CORE ;
  FOREIGN ao221_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 20.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 17.700 7.200 19.700 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.700 0.000 1.300 2.750 ;
        RECT 0.000 0.000 20.000 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 15.500 7.000 16.150 7.800 ;
        RECT 15.200 7.200 17.200 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.800 7.200 11.800 7.800 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 13.500 7.000 14.100 7.800 ;
        RECT 12.350 7.200 14.350 7.800 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.500 7.200 3.500 7.800 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 3.050 13.550 3.850 16.250 ;
        RECT 0.000 13.750 20.000 16.250 ;
        RECT 13.350 13.550 14.050 16.250 ;
        RECT 10.000 13.450 10.600 16.250 ;
        RECT 6.500 13.550 7.200 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.700 8.450 9.050 9.050 ;
    END
  END x
END ao221_4

MACRO ao221_3
  CLASS  CORE ;
  FOREIGN ao221_3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 18.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 7.200 2.250 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 3.050 0.000 3.650 2.750 ;
        RECT 0.000 0.000 18.750 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.050 7.200 5.050 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 16.500 7.200 18.500 7.800 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 14.050 5.950 16.050 6.550 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 11.050 7.200 13.050 7.800 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 4.350 13.550 5.050 16.250 ;
        RECT 0.000 13.750 18.750 16.250 ;
        RECT 12.500 13.550 13.200 16.250 ;
        RECT 7.750 13.550 8.450 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.100 7.200 10.150 7.800 ;
    END
  END x
END ao221_3

MACRO ao221_2
  CLASS  CORE ;
  FOREIGN ao221_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 17.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.650 7.200 2.650 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 17.500 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.250 7.200 5.250 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 15.250 7.200 17.250 7.800 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 13.400 6.250 14.000 7.800 ;
        RECT 13.400 7.200 14.750 7.800 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 10.700 7.200 12.700 7.800 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 4.350 13.550 5.050 16.250 ;
        RECT 0.000 13.750 17.500 16.250 ;
        RECT 7.750 13.550 8.450 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.100 8.450 10.150 9.050 ;
    END
  END x
END ao221_2

MACRO ao221_1
  CLASS  CORE ;
  FOREIGN ao221_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.800 8.450 4.800 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 15.000 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.300 8.450 2.300 9.050 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 12.650 7.200 14.650 7.800 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 11.450 9.700 13.450 10.300 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.900 7.200 11.900 7.800 ;
    END
  END e
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 3.800 13.550 4.500 16.250 ;
        RECT 0.000 13.750 15.000 16.250 ;
        RECT 7.200 13.550 7.900 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.550 8.450 9.600 9.050 ;
    END
  END x
END ao221_1

MACRO ao21_6
  CLASS  CORE ;
  FOREIGN ao21_6 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 20.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.500 4.600 10.100 5.300 ;
        RECT 9.050 4.700 11.250 5.300 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 6.650 0.000 7.250 3.550 ;
        RECT 0.000 0.000 20.000 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.900 4.700 3.900 5.300 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 16.000 8.450 18.250 9.050 ;
    END
  END c
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 9.200 13.450 9.900 16.250 ;
        RECT 0.000 13.750 20.000 16.250 ;
        RECT 12.600 13.450 13.300 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.450 8.450 11.600 9.050 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 14.350 7.200 19.350 7.800 ;
        RECT 14.350 7.200 14.950 10.350 ;
  END 
END ao21_6

MACRO ao21_5
  CLASS  CORE ;
  FOREIGN ao21_5 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 18.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.800 4.700 6.800 5.300 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 5.250 0.000 5.850 3.550 ;
        RECT 0.000 0.000 18.750 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.900 4.700 3.900 5.300 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 15.400 8.450 17.400 9.050 ;
    END
  END c
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 5.700 13.400 6.400 16.250 ;
        RECT 0.000 13.750 18.750 16.250 ;
        RECT 10.250 13.400 10.950 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.350 8.450 12.650 9.050 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 14.050 7.250 18.400 7.850 ;
        RECT 14.050 7.250 14.650 10.250 ;
        RECT 14.050 9.650 15.600 10.250 ;
  END 
END ao21_5

MACRO ao21_4
  CLASS  CORE ;
  FOREIGN ao21_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 16.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.900 4.700 5.900 5.300 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 4.600 0.000 5.200 3.550 ;
        RECT 0.000 0.000 16.250 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.050 4.700 3.050 5.300 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 13.000 7.200 15.000 7.800 ;
    END
  END c
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 5.800 13.450 6.500 16.250 ;
        RECT 0.000 13.750 16.250 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.200 4.700 11.750 5.300 ;
    END
  END x
END ao21_4

MACRO ao21_3
  CLASS  CORE ;
  FOREIGN ao21_3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.500 7.200 10.500 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 11.250 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.000 5.850 7.800 6.500 ;
        RECT 7.200 5.850 7.800 7.850 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.850 7.200 2.900 7.800 ;
    END
  END c
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 11.250 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.150 7.200 4.750 9.200 ;
        RECT 5.300 6.850 6.350 7.500 ;
        RECT 4.150 7.200 6.000 7.800 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 7.550 8.400 10.450 9.100 ;
  END 
END ao21_3

MACRO ao21_2
  CLASS  CORE ;
  FOREIGN ao21_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.350 10.950 0.950 11.650 ;
        RECT 0.350 10.950 2.350 11.550 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 6.350 0.000 6.950 2.700 ;
        RECT 0.000 0.000 10.000 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.100 9.700 3.100 10.300 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.450 5.950 4.450 6.550 ;
    END
  END c
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 10.000 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.250 8.450 9.600 9.050 ;
    END
  END x
END ao21_2

MACRO ao21_1
  CLASS  CORE ;
  FOREIGN ao21_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.400 5.950 4.750 6.550 ;
        RECT 4.150 7.300 4.950 7.900 ;
        RECT 4.150 5.950 4.750 7.900 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 7.500 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.200 7.250 2.800 9.150 ;
        RECT 2.200 7.250 3.650 7.850 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.350 5.950 2.350 6.550 ;
        RECT 1.550 5.950 2.350 6.600 ;
    END
  END c
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 7.500 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.750 5.950 7.150 6.550 ;
        RECT 6.550 5.950 7.150 9.100 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 3.550 8.500 6.050 9.100 ;
  END 
END ao21_1

MACRO ao211_5
  CLASS  CORE ;
  FOREIGN ao211_5 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 22.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.700 7.200 5.750 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 22.500 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.000 7.200 3.000 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 15.950 7.200 17.950 7.800 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 19.550 7.200 21.550 7.800 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 2.150 13.500 2.850 16.250 ;
        RECT 0.000 13.750 22.500 16.250 ;
        RECT 8.950 13.500 9.650 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.250 9.700 14.750 10.300 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 0.450 9.650 4.550 10.350 ;
  END 
END ao211_5

MACRO ao211_4
  CLASS  CORE ;
  FOREIGN ao211_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 20.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.700 7.200 5.700 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 20.000 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.500 7.200 2.850 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 15.500 8.450 17.500 9.050 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 17.150 7.200 19.150 7.800 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 20.000 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.100 8.450 14.750 9.050 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 9.500 7.200 16.100 7.800 ;
  END 
END ao211_4

MACRO ao211_3
  CLASS  CORE ;
  FOREIGN ao211_3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 17.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.650 7.200 5.700 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 17.500 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.850 7.200 2.850 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 11.900 7.200 13.900 7.800 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 14.900 7.200 17.000 7.800 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 17.500 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.550 8.450 10.700 9.050 ;
    END
  END x
END ao211_3

MACRO ao211_2
  CLASS  CORE ;
  FOREIGN ao211_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.100 5.950 10.100 6.550 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 15.000 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 10.950 5.900 11.550 7.900 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 12.450 5.950 14.450 6.550 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.850 7.200 2.850 7.800 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 15.000 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.950 7.200 4.600 7.900 ;
        RECT 3.950 7.200 7.350 7.800 ;
    END
  END x
END ao211_2

MACRO ao211_1
  CLASS  CORE ;
  FOREIGN ao211_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 10.050 7.250 10.650 9.050 ;
        RECT 9.400 8.450 10.650 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 13.750 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 11.300 7.200 13.300 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.350 7.200 4.350 7.800 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.350 7.100 1.850 7.900 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 13.750 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.850 7.200 8.750 7.800 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 1.550 8.450 6.450 9.050 ;
  END 
END ao211_1

MACRO and4i_5
  CLASS  CORE ;
  FOREIGN and4i_5 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 16.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.800 4.700 8.400 5.450 ;
        RECT 14.050 5.950 15.400 6.550 ;
        RECT 14.050 4.700 14.650 6.550 ;
        RECT 7.800 4.700 14.650 5.300 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 16.250 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.850 7.050 3.450 7.800 ;
        RECT 1.400 7.200 3.450 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.450 5.850 1.050 6.550 ;
        RECT 4.150 5.950 4.950 6.900 ;
        RECT 0.450 5.950 4.950 6.550 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.400 7.200 7.400 7.800 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 16.250 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 12.750 5.950 13.350 9.050 ;
        RECT 15.050 8.450 15.650 9.150 ;
        RECT 9.850 8.450 15.650 9.050 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 2.150 4.700 6.550 5.300 ;
        RECT 5.950 4.700 6.550 6.550 ;
        RECT 5.950 5.950 9.350 6.550 ;
        RECT 8.750 5.950 9.350 9.050 ;
        RECT 2.150 8.450 9.350 9.050 ;
  END 
END and4i_5

MACRO and4i_4
  CLASS  CORE ;
  FOREIGN and4i_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 10.000 6.600 10.950 7.800 ;
        RECT 10.000 7.200 11.750 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 13.750 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.600 7.200 2.600 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.450 5.400 1.050 6.550 ;
        RECT 0.450 5.950 4.150 6.550 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.900 7.200 6.000 7.800 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 13.750 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.150 8.450 12.750 9.050 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 2.150 4.700 7.650 5.300 ;
        RECT 7.050 4.700 7.650 10.300 ;
        RECT 0.450 9.700 7.650 10.300 ;
  END 
END and4i_4

MACRO and4i_3
  CLASS  CORE ;
  FOREIGN and4i_3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.400 8.450 11.650 9.100 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 5.350 0.000 5.950 2.800 ;
        RECT 0.000 0.000 12.500 2.500 ;
        RECT 6.650 0.000 7.250 2.800 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.850 5.950 2.950 6.550 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.550 7.200 4.550 7.800 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.600 5.950 6.650 6.550 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 12.500 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.300 7.200 10.450 7.800 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 5.150 7.200 7.750 7.800 ;
        RECT 5.150 7.200 5.750 9.050 ;
        RECT 0.450 8.450 5.750 9.050 ;
  END 
END and4i_3

MACRO and4i_2
  CLASS  CORE ;
  FOREIGN and4i_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.750 5.700 5.850 6.300 ;
        RECT 5.300 5.950 6.550 6.550 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 10.000 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 5.850 1.750 6.650 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.350 8.450 9.650 9.050 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.450 4.900 4.050 6.900 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 1.000 13.500 1.600 16.250 ;
        RECT 0.000 13.750 10.000 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.850 3.450 7.800 4.050 ;
        RECT 7.200 5.950 9.150 6.550 ;
        RECT 7.200 3.450 7.800 6.550 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 0.350 3.450 2.850 4.050 ;
        RECT 2.250 3.800 5.350 4.400 ;
        RECT 4.750 3.800 5.350 5.200 ;
        RECT 4.750 4.600 6.450 5.200 ;
        RECT 2.250 3.450 2.850 6.650 ;
  END 
END and4i_2

MACRO and4i_1
  CLASS  CORE ;
  FOREIGN and4i_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.250 8.450 6.250 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 3.850 0.000 4.450 2.800 ;
        RECT 0.000 0.000 8.750 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.400 8.450 2.400 9.050 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.050 5.950 3.050 6.550 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.800 4.700 4.800 5.300 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 1.200 13.550 1.900 16.250 ;
        RECT 0.000 13.750 8.750 16.250 ;
        RECT 4.750 13.450 5.350 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.550 5.950 8.300 6.550 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 0.350 7.150 6.850 7.750 ;
        RECT 0.350 7.150 3.550 7.800 ;
        RECT 2.950 7.150 3.550 9.000 ;
  END 
END and4i_1

MACRO and4_5
  CLASS  CORE ;
  FOREIGN and4_5 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.900 8.450 11.650 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 3.650 0.000 4.250 2.800 ;
        RECT 0.000 0.000 12.500 2.500 ;
        RECT 5.250 0.000 5.850 2.800 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.150 7.200 10.300 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.550 7.300 7.200 9.050 ;
        RECT 5.850 8.450 7.200 9.050 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.400 7.200 5.400 7.800 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 12.500 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 7.200 2.750 7.800 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 0.850 9.700 12.150 10.300 ;
  END 
END and4_5

MACRO and4_4
  CLASS  CORE ;
  FOREIGN and4_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.400 7.200 5.400 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 11.250 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.950 8.350 6.600 9.050 ;
        RECT 5.350 8.450 7.350 9.050 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.100 7.200 9.400 7.800 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.900 8.450 10.900 9.050 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 6.950 13.500 7.550 16.250 ;
        RECT 0.000 13.750 11.250 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.450 7.200 2.750 7.800 ;
    END
  END x
END and4_4

MACRO and4_3
  CLASS  CORE ;
  FOREIGN and4_3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.200 8.450 4.200 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 10.000 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.350 5.950 6.350 6.550 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.250 8.450 7.250 9.050 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.750 8.450 9.750 9.050 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 2.150 13.100 2.750 16.250 ;
        RECT 0.000 13.750 10.000 16.250 ;
        RECT 5.550 13.100 6.150 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.450 5.950 2.450 6.550 ;
    END
  END x
END and4_3

MACRO and4_2
  CLASS  CORE ;
  FOREIGN and4_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.500 7.200 6.750 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 8.750 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.400 5.950 4.000 7.250 ;
        RECT 3.400 5.950 6.400 6.550 ;
        RECT 3.000 6.650 4.000 7.250 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.100 8.450 3.100 9.050 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 5.950 2.250 6.550 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 8.750 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.350 9.700 8.350 10.300 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 6.500 8.400 7.100 9.050 ;
        RECT 4.100 8.450 7.100 9.050 ;
  END 
END and4_2

MACRO and4_1
  CLASS  CORE ;
  FOREIGN and4_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.700 5.950 5.800 6.550 ;
        RECT 5.200 5.950 5.800 7.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 8.750 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.050 8.450 3.750 9.050 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.850 7.200 4.400 7.800 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.350 4.700 4.800 5.300 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 8.750 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.400 7.200 8.400 7.800 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 4.250 8.450 7.150 9.050 ;
  END 
END and4_1

MACRO and3i_5
  CLASS  CORE ;
  FOREIGN and3i_5 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.900 7.200 8.400 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 15.000 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 10.850 7.200 12.900 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.400 4.700 9.100 5.400 ;
        RECT 12.150 4.700 12.800 5.400 ;
        RECT 8.400 4.700 12.800 5.300 ;
    END
  END c
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 15.000 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.450 4.700 1.100 5.400 ;
        RECT 0.450 4.700 6.650 5.300 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 1.750 5.950 14.300 6.550 ;
  END 
END and3i_5

MACRO and3i_4
  CLASS  CORE ;
  FOREIGN and3i_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.600 7.200 3.600 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 12.500 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 10.250 8.450 12.250 9.050 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.300 4.700 12.150 5.300 ;
    END
  END c
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 12.500 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.350 9.700 6.250 10.300 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 6.200 3.400 9.550 4.000 ;
        RECT 6.200 3.400 6.800 5.400 ;
        RECT 6.750 7.150 10.350 7.750 ;
        RECT 6.750 7.150 7.350 9.050 ;
        RECT 1.100 8.450 7.350 9.050 ;
  END 
END and3i_4

MACRO and3i_3
  CLASS  CORE ;
  FOREIGN and3i_3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.150 4.700 2.100 6.550 ;
        RECT 4.750 5.900 5.450 6.650 ;
        RECT 4.750 4.700 5.350 6.650 ;
        RECT 1.150 4.700 5.350 5.300 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 10.000 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.750 6.700 8.350 7.800 ;
        RECT 7.750 7.200 9.600 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.400 4.700 7.100 6.550 ;
        RECT 6.400 4.700 8.000 5.300 ;
    END
  END c
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 10.000 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.950 7.200 1.650 10.250 ;
        RECT 0.950 7.200 3.950 7.800 ;
        RECT 3.350 5.900 3.950 7.800 ;
        RECT 0.950 9.600 3.700 10.250 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 2.250 8.300 2.850 9.050 ;
        RECT 2.250 8.450 9.650 9.050 ;
  END 
END and3i_3

MACRO and3i_2
  CLASS  CORE ;
  FOREIGN and3i_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.350 4.700 5.350 5.300 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 10.000 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.150 4.700 9.150 5.300 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.500 5.950 7.500 6.550 ;
    END
  END c
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 10.000 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.850 5.950 3.950 6.550 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 3.100 7.050 3.800 7.800 ;
        RECT 3.100 7.200 9.400 7.800 ;
  END 
END and3i_2

MACRO and3i_1
  CLASS  CORE ;
  FOREIGN and3i_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.900 8.450 2.900 9.050 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 7.500 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.750 7.200 6.750 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.250 5.950 5.250 6.550 ;
    END
  END c
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 7.500 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.400 5.950 2.750 6.550 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 4.700 8.450 7.150 9.050 ;
  END 
END and3i_1

MACRO and3_5
  CLASS  CORE ;
  FOREIGN and3_5 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.700 5.950 9.700 6.550 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 10.000 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.700 7.200 7.700 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.350 5.950 4.950 6.550 ;
        RECT 4.150 5.950 4.950 7.150 ;
    END
  END c
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 10.000 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.600 7.200 2.600 7.800 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 3.250 8.000 3.900 9.200 ;
        RECT 3.250 8.600 9.650 9.200 ;
  END 
END and3_5

MACRO and3_4
  CLASS  CORE ;
  FOREIGN and3_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.750 7.200 9.750 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 10.000 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.850 5.950 7.850 6.550 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.350 7.200 5.350 7.800 ;
    END
  END c
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 10.000 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.850 5.950 3.300 6.550 ;
    END
  END x
END and3_4

MACRO and3_3
  CLASS  CORE ;
  FOREIGN and3_3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.500 5.950 7.200 6.600 ;
        RECT 6.500 5.950 8.500 6.550 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 8.750 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.500 7.200 6.500 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.150 5.950 4.200 6.550 ;
        RECT 3.550 5.950 4.200 6.600 ;
    END
  END c
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 2.550 13.600 3.250 16.250 ;
        RECT 0.000 13.750 8.750 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.350 8.500 0.950 10.300 ;
        RECT 0.350 9.700 1.850 10.300 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 1.650 8.450 8.400 9.050 ;
  END 
END and3_3

MACRO and3_2
  CLASS  CORE ;
  FOREIGN and3_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.000 7.200 8.000 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 8.750 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.500 7.200 5.500 7.800 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.550 9.700 4.550 10.300 ;
    END
  END c
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 8.750 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 7.200 2.250 7.800 ;
    END
  END x
END and3_2

MACRO and3_1
  CLASS  CORE ;
  FOREIGN and3_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.150 5.950 7.150 6.550 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 7.500 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.200 8.450 6.250 9.050 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.600 5.950 4.600 6.550 ;
    END
  END c
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 5.700 13.450 6.400 16.250 ;
        RECT 0.000 13.750 7.500 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 8.450 2.250 9.050 ;
    END
  END x
END and3_1

MACRO and2_8
  CLASS  CORE ;
  FOREIGN and2_8 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.600 5.950 11.750 6.550 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 6.250 0.000 6.950 2.600 ;
        RECT 0.000 0.000 12.500 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.950 4.650 7.200 5.500 ;
        RECT 5.950 4.650 11.400 5.250 ;
    END
  END b
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 12.500 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.750 4.700 4.850 5.300 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 1.800 7.200 11.650 7.800 ;
  END 
END and2_8

MACRO and2_6
  CLASS  CORE ;
  FOREIGN and2_6 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.000 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.500 5.950 7.100 6.650 ;
        RECT 6.500 5.950 8.500 6.550 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 10.000 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.800 5.950 5.400 6.650 ;
        RECT 4.000 5.950 6.000 6.550 ;
    END
  END b
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 10.000 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.850 5.950 3.350 6.550 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 0.850 8.450 9.600 9.050 ;
  END 
END and2_6

MACRO and2_5
  CLASS  CORE ;
  FOREIGN and2_5 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.400 5.950 8.400 6.550 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 8.750 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.900 5.950 5.900 6.550 ;
    END
  END b
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 8.750 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.400 5.950 3.400 6.550 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 1.000 8.450 8.300 9.050 ;
  END 
END and2_5

MACRO and2_4
  CLASS  CORE ;
  FOREIGN and2_4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.000 5.950 8.000 6.550 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 8.750 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.500 5.950 5.500 6.550 ;
    END
  END b
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 8.750 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.000 5.950 3.000 6.550 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 3.350 8.300 4.050 9.050 ;
        RECT 3.350 8.450 8.400 9.050 ;
  END 
END and2_4

MACRO and2_3
  CLASS  CORE ;
  FOREIGN and2_3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.050 7.200 7.050 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 7.500 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.350 7.200 4.350 7.800 ;
    END
  END b
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 7.500 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 9.700 2.250 10.300 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 2.750 9.700 6.800 10.300 ;
        RECT 1.650 8.450 7.150 9.050 ;
  END 
END and2_3

MACRO and2_2
  CLASS  CORE ;
  FOREIGN and2_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.850 7.200 5.850 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 7.500 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.300 9.700 5.300 10.300 ;
    END
  END b
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 7.500 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 7.200 2.250 7.800 ;
    END
  END x
END and2_2

MACRO and2_1
  CLASS  CORE ;
  FOREIGN and2_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.400 4.700 5.450 5.300 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 6.250 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.150 7.200 4.150 7.800 ;
    END
  END b
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 6.250 16.250 ;
    END
  END vdd!
  PIN x
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.550 4.700 2.550 5.300 ;
    END
  END x
  OBS 
      LAYER Metal1 ;
        RECT 2.000 8.450 4.800 9.050 ;
  END 
END and2_1

MACRO adhalf_2
  CLASS  CORE ;
  FOREIGN adhalf_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 17.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.700 5.950 2.700 6.550 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 17.500 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.000 5.950 11.000 6.550 ;
    END
  END b
  PIN s
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 13.150 5.850 14.050 6.600 ;
        RECT 13.450 7.800 14.150 8.650 ;
        RECT 13.450 5.850 14.050 8.650 ;
    END
  END s
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 17.500 16.250 ;
    END
  END vdd!
  PIN co
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.550 5.350 6.150 6.550 ;
        RECT 5.550 5.950 7.850 6.550 ;
    END
  END co
  OBS 
      LAYER Metal1 ;
        RECT 4.300 5.950 4.900 8.300 ;
        RECT 4.300 7.700 9.050 8.300 ;
        RECT 15.500 8.300 16.100 9.750 ;
        RECT 11.850 9.150 16.100 9.750 ;
  END 
END adhalf_2

MACRO adhalf_1
  CLASS  CORE ;
  FOREIGN adhalf_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.450 7.750 9.050 10.400 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 12.500 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.350 8.450 5.450 9.050 ;
    END
  END b
  PIN s
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.450 7.200 6.600 7.800 ;
        RECT 5.450 9.700 6.600 10.300 ;
        RECT 6.000 7.200 6.600 10.300 ;
    END
  END s
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 13.750 12.500 16.250 ;
    END
  END vdd!
  PIN co
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 10.550 7.250 11.150 10.300 ;
        RECT 10.550 9.700 12.050 10.300 ;
    END
  END co
  OBS 
      LAYER Metal1 ;
        RECT 0.250 6.300 0.950 6.900 ;
        RECT 0.250 6.300 0.850 10.150 ;
        RECT 0.250 9.550 1.050 10.150 ;
        RECT 2.450 6.100 12.250 6.700 ;
        RECT 2.450 6.100 3.050 7.800 ;
        RECT 11.650 6.100 12.250 8.950 ;
  END 
END adhalf_1

MACRO adfullm_2
  CLASS  CORE ;
  FOREIGN adfullm_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 27.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 3.400 2.050 4.100 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 9.500 0.000 10.100 2.700 ;
        RECT 0.000 0.000 27.500 2.500 ;
        RECT 12.850 0.000 13.450 2.700 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.050 7.200 11.050 7.800 ;
    END
  END b
  PIN s
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 21.450 4.550 22.900 5.150 ;
        RECT 21.750 8.450 22.900 9.050 ;
        RECT 22.300 4.550 22.900 9.050 ;
    END
  END s
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 9.500 13.550 10.100 16.250 ;
        RECT 0.000 13.750 27.500 16.250 ;
    END
  END vdd!
  PIN ci
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 24.650 7.200 26.650 7.800 ;
    END
  END ci
  PIN co
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 13.850 6.050 14.450 9.050 ;
        RECT 13.850 8.350 16.050 9.050 ;
        RECT 13.850 6.050 15.150 6.650 ;
    END
  END co
  OBS 
      LAYER Metal1 ;
        RECT 3.300 7.500 6.100 8.100 ;
        RECT 6.100 6.400 7.200 7.000 ;
        RECT 6.600 6.400 7.200 9.200 ;
        RECT 6.100 8.600 7.200 9.200 ;
        RECT 3.300 3.100 7.850 3.700 ;
        RECT 3.300 3.100 3.900 5.900 ;
        RECT 1.000 5.300 3.900 5.900 ;
        RECT 4.400 4.200 11.800 4.800 ;
        RECT 14.950 3.000 15.550 4.450 ;
        RECT 12.750 3.850 15.550 4.450 ;
        RECT 5.000 5.300 13.350 5.900 ;
        RECT 5.000 5.300 5.600 7.000 ;
        RECT 2.200 6.400 5.600 7.000 ;
        RECT 12.750 3.850 13.350 7.800 ;
        RECT 2.200 6.400 2.800 9.200 ;
        RECT 2.200 8.600 3.300 9.200 ;
        RECT 17.150 8.250 20.700 8.850 ;
        RECT 21.200 6.150 21.800 7.750 ;
        RECT 14.950 7.150 21.800 7.750 ;
        RECT 23.500 8.450 27.050 9.050 ;
        RECT 20.000 3.450 27.150 4.050 ;
        RECT 26.550 3.450 27.150 5.550 ;
        RECT 20.000 3.450 20.600 6.650 ;
        RECT 18.450 6.050 20.600 6.650 ;
  END 
END adfullm_2

MACRO adfullm_1
  CLASS  CORE ;
  FOREIGN adfullm_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 23.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.250 3.400 2.050 4.100 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 9.500 0.000 10.100 3.150 ;
        RECT 0.000 0.000 23.750 2.500 ;
        RECT 16.300 0.000 16.900 2.700 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.100 7.150 9.700 7.800 ;
        RECT 8.550 7.200 10.550 7.800 ;
    END
  END b
  PIN s
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 19.700 6.400 21.550 7.000 ;
        RECT 19.700 8.600 21.550 9.200 ;
        RECT 20.850 6.400 21.550 9.200 ;
    END
  END s
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 9.500 13.550 10.100 16.250 ;
        RECT 0.000 13.750 23.750 16.250 ;
        RECT 19.650 13.600 20.350 16.250 ;
        RECT 16.300 13.550 16.900 16.250 ;
    END
  END vdd!
  PIN ci
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 16.600 7.150 17.300 7.800 ;
        RECT 15.900 7.200 17.900 7.800 ;
    END
  END ci
  PIN co
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 12.200 6.400 12.900 9.200 ;
        RECT 12.200 8.600 13.500 9.200 ;
        RECT 12.200 6.400 13.500 7.000 ;
    END
  END co
  OBS 
      LAYER Metal1 ;
        RECT 3.300 7.500 6.100 8.100 ;
        RECT 6.100 6.400 7.200 7.000 ;
        RECT 6.600 6.400 7.200 9.200 ;
        RECT 6.100 8.600 7.200 9.200 ;
        RECT 3.300 3.100 7.850 3.700 ;
        RECT 3.300 3.100 3.900 5.900 ;
        RECT 1.000 5.300 3.900 5.900 ;
        RECT 4.400 4.200 11.800 4.800 ;
        RECT 14.750 6.000 19.000 6.600 ;
        RECT 18.400 6.000 19.000 8.100 ;
        RECT 14.750 6.000 15.350 8.100 ;
        RECT 13.500 7.500 15.350 8.100 ;
        RECT 18.400 7.500 19.700 8.100 ;
        RECT 14.600 4.900 22.000 5.500 ;
        RECT 19.150 3.250 19.750 4.400 ;
        RECT 13.450 3.800 23.300 4.400 ;
        RECT 13.450 3.250 14.050 5.900 ;
        RECT 5.000 5.300 14.050 5.900 ;
        RECT 5.000 5.300 5.600 7.000 ;
        RECT 2.200 6.400 5.600 7.000 ;
        RECT 22.700 3.800 23.300 7.800 ;
        RECT 2.200 6.400 2.800 9.200 ;
        RECT 2.200 8.600 3.300 9.200 ;
  END 
END adfullm_1

MACRO adfull_2
  CLASS  CORE ;
  FOREIGN adfull_2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 28.750 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.750 7.200 2.800 7.800 ;
        RECT 2.200 6.600 11.900 7.200 ;
        RECT 4.050 6.350 4.700 7.200 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 19.200 0.000 19.800 2.700 ;
        RECT 0.000 0.000 28.750 2.500 ;
        RECT 26.000 0.000 26.600 2.700 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.350 7.700 6.950 9.050 ;
        RECT 3.150 8.450 6.950 9.050 ;
    END
  END b
  PIN s
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 15.800 6.750 16.400 9.050 ;
        RECT 15.800 8.450 16.850 9.050 ;
    END
  END s
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 7.300 13.550 7.900 16.250 ;
        RECT 0.000 13.750 28.750 16.250 ;
        RECT 26.000 13.550 26.600 16.250 ;
        RECT 10.700 13.550 11.300 16.250 ;
    END
  END vdd!
  PIN ci
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 25.800 7.100 27.300 7.900 ;
    END
  END ci
  PIN co
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 22.100 6.150 22.700 9.050 ;
        RECT 22.100 8.450 23.200 9.050 ;
        RECT 22.100 6.150 23.200 6.750 ;
    END
  END co
  OBS 
      LAYER Metal1 ;
        RECT 0.350 8.450 2.650 9.050 ;
        RECT 9.000 8.450 13.000 9.050 ;
        RECT 9.400 4.400 19.400 5.000 ;
        RECT 18.800 4.400 19.400 6.600 ;
        RECT 4.750 4.400 8.900 5.000 ;
        RECT 8.300 4.400 8.900 6.100 ;
        RECT 8.300 5.500 18.100 6.100 ;
        RECT 17.500 5.500 18.100 7.700 ;
        RECT 17.500 7.100 20.500 7.700 ;
        RECT 20.900 4.850 21.600 5.500 ;
        RECT 21.000 4.850 21.600 8.850 ;
        RECT 20.900 8.250 21.600 8.850 ;
        RECT 0.350 3.300 23.100 3.900 ;
        RECT 0.350 3.300 0.950 4.650 ;
        RECT 22.500 3.300 23.100 5.500 ;
        RECT 22.500 4.900 26.200 5.500 ;
        RECT 25.600 4.900 26.200 6.600 ;
        RECT 23.200 7.250 25.050 7.850 ;
        RECT 24.450 7.250 25.050 9.000 ;
        RECT 27.800 6.950 28.400 9.000 ;
        RECT 24.450 8.400 28.400 9.000 ;
  END 
END adfull_2

MACRO adfull_1
  CLASS  CORE ;
  FOREIGN adfull_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 26.250 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.450 6.650 9.050 7.800 ;
        RECT 1.900 7.200 9.050 7.800 ;
    END
  END a
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 26.250 2.500 ;
    END
  END vss!
  PIN b
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.800 7.150 10.400 9.050 ;
        RECT 3.150 8.450 10.400 9.050 ;
    END
  END b
  PIN s
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 14.300 6.750 14.900 9.050 ;
        RECT 14.300 8.450 15.500 9.050 ;
    END
  END s
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 9.200 13.550 9.800 16.250 ;
        RECT 0.000 13.750 26.250 16.250 ;
    END
  END vdd!
  PIN ci
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 24.000 8.450 26.000 9.050 ;
    END
  END ci
  PIN co
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 21.200 6.650 21.800 9.050 ;
        RECT 20.700 8.450 21.800 9.050 ;
    END
  END co
  OBS 
      LAYER Metal1 ;
        RECT 0.350 8.450 2.650 9.050 ;
        RECT 8.300 4.450 17.900 5.050 ;
        RECT 17.300 4.450 17.900 7.400 ;
        RECT 5.300 4.700 7.800 5.300 ;
        RECT 7.200 4.700 7.800 6.150 ;
        RECT 7.200 5.550 16.600 6.150 ;
        RECT 16.000 5.550 16.600 8.500 ;
        RECT 16.000 7.900 19.000 8.500 ;
        RECT 19.500 6.400 20.100 9.100 ;
        RECT 1.150 3.350 24.800 3.950 ;
        RECT 1.150 3.350 1.750 4.750 ;
        RECT 24.200 3.350 24.800 7.800 ;
  END 
END adfull_1

MACRO sdffn_1
  CLASS  CORE ;
  FOREIGN sdffn_1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 22.500 BY 16.250 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 20.150 5.950 22.150 6.550 ;
    END
  END q
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 3.100 0.000 3.700 2.650 ;
        RECT 0.000 0.000 22.500 2.500 ;
        RECT 19.800 0.000 20.400 2.700 ;
        RECT 13.700 0.000 14.300 2.600 ;
        RECT 11.450 0.000 12.050 2.600 ;
    END
  END vss!
  PIN ckb
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.650 3.450 13.350 4.050 ;
    END
  END ckb
  PIN se
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.050 6.650 4.050 7.250 ;
        RECT 3.450 8.550 4.100 9.150 ;
        RECT 3.450 5.950 4.050 9.150 ;
    END
  END se
  PIN d
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.100 6.900 5.700 9.050 ;
        RECT 4.700 8.450 5.700 9.050 ;
    END
  END d
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 3.450 13.550 4.050 16.250 ;
        RECT 0.000 13.750 22.500 16.250 ;
        RECT 19.750 13.550 20.350 16.250 ;
        RECT 11.800 13.550 12.400 16.250 ;
    END
  END vdd!
  PIN qb
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 19.500 8.450 21.500 9.050 ;
    END
  END qb
  PIN sdi
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.500 7.500 2.100 9.050 ;
        RECT 1.500 8.450 2.900 9.050 ;
    END
  END sdi
  OBS 
      LAYER Metal1 ;
        RECT 0.350 5.950 0.950 10.300 ;
        RECT 6.200 5.950 6.800 10.300 ;
        RECT 0.350 9.700 6.800 10.300 ;
        RECT 7.300 5.950 8.950 6.550 ;
        RECT 7.300 5.950 7.900 10.300 ;
        RECT 7.300 9.700 8.900 10.300 ;
        RECT 9.150 8.400 9.800 9.050 ;
        RECT 9.150 8.450 17.750 9.050 ;
        RECT 8.400 7.050 10.900 7.650 ;
        RECT 15.600 7.150 18.400 7.750 ;
        RECT 10.250 7.350 16.200 7.950 ;
  END 
END sdffn_1

#END LIBRARY
#******
# Preview export LEF
#
#	 Preview sub-version 4.4.3.100.44
#
# TECH LIB NAME: cdr3_dev
# TECH FILE NAME: techfile.cds
#******
# metal 5 update was done for all corner cells, fill cells
#         allvdd,allvss,outvss,outvdd and for inbuf3_16 and
#         iobuf3_16_12 cells others were not !! be changed
#         u.j. march 2002
#         iobuf3_16_8 / iobuf3_16pu_8        port  CLASS CORE;
#         iobuf2_16_12 / inbuf2_16           port  CLASS CORE;
#         iobuf3_16_12 / iobuf3_16pu_12      port  CLASS CORE;
#         inbuf3_16pu
#         inbufs3_16pu

MACRO allvdd
    CLASS PAD ;
    FOREIGN allvdd  0.00 -38.75 N  ;
    ORIGIN 0.00 39.15 ;
    SIZE 115.00 BY 600.00 ;
    SYMMETRY x y r90 ;
    SITE io_site ;
    PIN pad USE POWER ; DIRECTION INPUT ;
        PORT
        LAYER Metal5 ;
        RECT  3.00 383.00 112.00 544.25 ;
        END
    END pad
    OBS
        LAYER Metal1 ;
        RECT  0.25 -0.40 114.75 560.00 ;
        LAYER Metal2 ;
        RECT  0.33 0.33 114.68 559.92 ;
        LAYER Metal3 ;
        RECT  0.33 0.33 114.68 559.92 ;
        LAYER Metal4 ;
        RECT  0.33 0.33 114.68 559.92 ;
        LAYER Metal5 ;
        RECT  0.33 0.33 114.68 559.92 ;
    END
END allvdd

MACRO allvss
    CLASS PAD ;
    FOREIGN allvss  0.00 -38.75 N  ;
    ORIGIN 0.00 39.15 ;
    SIZE 115.00 BY 600.00 ;
    SYMMETRY x y r90 ;
    SITE io_site ;
    PIN pad USE power ; DIRECTION INPUT ;
        PORT
        LAYER Metal5 ;
        RECT  3.00 383.00 112.00 544.25 ;
        END
    END pad
    OBS
        LAYER Metal1 ;
        RECT  0.25 -0.40 114.75 560.00 ;
        LAYER Metal2 ;
        RECT  0.33 0.33 114.68 559.92 ;
        LAYER Metal3 ;
        RECT  0.33 0.33 114.68 559.92 ;
        LAYER Metal4 ;
        RECT  0.33 0.33 114.68 559.92 ;
        LAYER Metal5 ;
        RECT  0.33 0.33 114.68 559.92 ;
    END
END allvss







MACRO inbuf2_16
    CLASS PAD ;
    FOREIGN inbuf2_16  0.00 -38.75 N  ;
    ORIGIN 0.00 39.15 ;
    SIZE 115.00 BY 600.00 ;
    SYMMETRY x y r90 ;
    SITE io_site ;
    PIN di  USE SIGNAL ; DIRECTION OUTPUT ;
        PORT
        LAYER Metal1 ;
        RECT  87.15 -0.40 87.75 0.30 ;
        END
    END di
    PIN pad USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal3 ;
        RECT  3.00 383.00 112.00 544.25 ;
        END
    END pad
    PIN vdd!
        USE power ;  DIRECTION INOUT ;
        PORT
        CLASS CORE ;
        LAYER Metal2 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        LAYER Metal3 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        END
    END vdd!
    PIN vss!
        USE ground ;  DIRECTION INOUT ;
        PORT
        CLASS CORE ;
        LAYER Metal2 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        LAYER Metal3 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        END
    END vss!

    OBS
        LAYER Metal1 ;
        RECT  88.35 -0.40 114.75 560.00 ;
        RECT  86.55 0.90 88.35 560.00 ;
        RECT  0.25 -0.40 86.55 560.00 ;
        LAYER Metal2 ;
        RECT  0.33 0.33 114.68 559.92 ;
        LAYER Metal3 ;
        RECT  114.65 0.33 114.68 559.92 ;
        RECT  103.70 2.20 114.65 559.92 ;
        RECT  0.33 0.33 2.20 0.60 ;
        RECT  0.33 54.65 2.20 59.75 ;
        RECT  0.33 108.90 2.20 109.60 ;
        RECT  0.33 241.90 2.20 242.60 ;
        RECT  0.33 380.90 2.20 559.92 ;
        RECT  2.20 0.33 103.70 559.92 ;
    END
END inbuf2_16

MACRO inbuf2_16pd
    CLASS PAD ;
    FOREIGN inbuf2_16pd  0.00 -38.75 N  ;
    ORIGIN 0.00 39.15 ;
    SIZE 115.00 BY 600.00 ;
    SYMMETRY x y r90 ;
    SITE io_site ;
    PIN di  USE SIGNAL ; DIRECTION OUTPUT ;
        PORT
        LAYER Metal1 ;
        RECT  87.15 -0.40 87.75 0.30 ;
        END
    END di
    PIN pad USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal3 ;
        RECT  3.00 383.00 112.00 544.25 ;
        END
    END pad
    PIN vdd!
        USE power ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        LAYER Metal3 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        END
    END vdd!
    PIN vss!
        USE ground ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        LAYER Metal3 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        END
    END vss!
    OBS
        LAYER Metal1 ;
        RECT  88.35 -0.40 114.75 560.00 ;
        RECT  86.55 0.90 88.35 560.00 ;
        RECT  0.25 -0.40 86.55 560.00 ;
        LAYER Metal2 ;
        RECT  0.33 0.33 114.68 559.92 ;
        LAYER Metal3 ;
        RECT  114.65 0.33 114.68 559.92 ;
        RECT  103.70 2.20 114.65 559.92 ;
        RECT  4.05 2.20 14.70 559.92 ;
        RECT  2.20 0.33 4.05 559.92 ;
        RECT  0.33 0.33 2.20 59.75 ;
        RECT  0.33 108.90 2.20 109.60 ;
        RECT  0.33 241.90 2.20 242.60 ;
        RECT  0.33 380.90 2.20 559.92 ;
        RECT  14.70 0.33 103.70 559.92 ;
    END
END inbuf2_16pd

MACRO inbuf2_16pu
    CLASS PAD ;
    FOREIGN inbuf2_16pu  0.00 -38.75 N  ;
    ORIGIN 0.00 39.15 ;
    SIZE 115.00 BY 600.00 ;
    SYMMETRY x y r90 ;
    SITE io_site ;
    PIN di  USE SIGNAL ; DIRECTION OUTPUT ;
        PORT
        LAYER Metal1 ;
        RECT  87.15 -0.40 87.75 0.30 ;
        END
    END di
    PIN pad USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal3 ;
        RECT  3.00 383.00 112.00 544.25 ;
        END
    END pad
    PIN vdd!
        USE power ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        LAYER Metal3 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        END
    END vdd!
    PIN vss!
        USE ground ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        LAYER Metal3 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        END
    END vss!
    OBS
        LAYER Metal1 ;
        RECT  88.35 -0.40 114.75 560.00 ;
        RECT  86.55 0.90 88.35 560.00 ;
        RECT  0.25 -0.40 86.55 560.00 ;
        LAYER Metal2 ;
        RECT  0.33 0.33 114.68 559.92 ;
        LAYER Metal3 ;
        RECT  114.65 0.33 114.68 559.92 ;
        RECT  103.70 2.20 114.65 559.92 ;
        RECT  4.05 2.20 14.70 559.92 ;
        RECT  2.20 0.33 4.05 559.92 ;
        RECT  0.33 0.33 2.20 59.75 ;
        RECT  0.33 108.90 2.20 109.60 ;
        RECT  0.33 241.90 2.20 242.60 ;
        RECT  0.33 380.90 2.20 559.92 ;
        RECT  14.70 0.33 103.70 559.92 ;
    END
END inbuf2_16pu



MACRO inbuf3_16
    CLASS PAD ;
    FOREIGN inbuf3_16  0.00 -38.75 N  ;
    ORIGIN 0.00 39.15 ;
    SIZE 115.00 BY 600.00 ;
    SYMMETRY x y r90 ;
    SITE io_site ;
    PIN di  USE SIGNAL ; DIRECTION OUTPUT ;
        PORT
        LAYER Metal1 ;
        RECT  87.15 -0.40 87.75 0.30 ;
        END
    END di
    PIN pad USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal5 ;
        RECT  3.00 383.00 112.00 544.25 ;
        END
    END pad
    PIN vdd!
        USE power ;  DIRECTION INOUT ;
        PORT
        CLASS CORE ;
        LAYER Metal2 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        LAYER Metal3 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        END
    END vdd!
    PIN vss!
        USE ground ;  DIRECTION INOUT ;
        PORT
        CLASS CORE ;
        LAYER Metal2 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        LAYER Metal3 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        END
    END vss!
    OBS
        LAYER Metal1 ;
        RECT  88.35 -0.40 114.75 560.00 ;
        RECT  86.55 0.90 88.35 560.00 ;
        RECT  0.25 -0.40 86.55 560.00 ;
        LAYER Metal2 ;
        RECT  0.33 0.33 114.68 559.92 ;
        LAYER Metal3 ;
        RECT  114.65 0.33 114.68 559.92 ;
        RECT  103.70 2.20 114.65 559.92 ;
        RECT  4.05 2.20 14.70 559.92 ;
        RECT  2.20 0.33 4.05 559.92 ;
        RECT  0.33 0.33 2.20 59.75 ;
        RECT  0.33 108.90 2.20 109.60 ;
        RECT  0.33 241.90 2.20 242.60 ;
        RECT  0.33 380.90 2.20 559.92 ;
        RECT  14.70 0.33 103.70 559.92 ;
        LAYER Metal4 ;
        RECT  0.33 0.33 114.68 559.92 ;
        LAYER Metal5 ;
        RECT  114.65 0.33 114.68 559.92 ;
        RECT  103.70 2.20 114.65 559.92 ;
        RECT  4.05 2.20 14.70 559.92 ;
        RECT  2.20 0.33 4.05 559.92 ;
        RECT  0.33 0.33 2.20 59.75 ;
        RECT  0.33 108.90 2.20 109.60 ;
        RECT  0.33 241.90 2.20 242.60 ;
        RECT  0.33 380.90 2.20 559.92 ;
        RECT  14.70 0.33 103.70 559.92 ;

    END
END inbuf3_16


MACRO analog_gnd
    CLASS PAD ;
    FOREIGN analog_gnd  0.00 -38.75 N  ;
    ORIGIN 0.00 39.15 ;
    SIZE 115.00 BY 600.00 ;
    SYMMETRY x y r90 ;
    SITE io_site ;
    PIN gnda!
        USE ground ;  DIRECTION INOUT ;
        PORT
        CLASS CORE ;
        LAYER Metal1 ;
        RECT  14.00 -0.40 114.00 1.55 ;
        LAYER Metal2 ;
        RECT  14.00 -0.40 114.00 1.55 ;
        END
    END gnda!
    OBS
        LAYER Metal1 ;
        RECT  88.35 -0.40 114.75 560.00 ;
        RECT  86.55 0.90 88.35 560.00 ;
        RECT  0.25 -0.40 86.55 560.00 ;
        LAYER Metal2 ;
        RECT  0.33 0.33 114.68 559.92 ;
        LAYER Metal3 ;
        RECT  114.65 0.33 114.68 559.92 ;
        RECT  103.70 2.20 114.65 559.92 ;
        RECT  4.05 2.20 14.70 559.92 ;
        RECT  2.20 0.33 4.05 559.92 ;
        RECT  0.33 0.33 2.20 59.75 ;
        RECT  0.33 108.90 2.20 109.60 ;
        RECT  0.33 241.90 2.20 242.60 ;
        RECT  0.33 380.90 2.20 559.92 ;
        RECT  14.70 0.33 103.70 559.92 ;
        LAYER Metal4 ;
        RECT  0.33 0.33 114.68 559.92 ;
        LAYER Metal5 ;
        RECT  114.65 0.33 114.68 559.92 ;
        RECT  103.70 2.20 114.65 559.92 ;
        RECT  4.05 2.20 14.70 559.92 ;
        RECT  2.20 0.33 4.05 559.92 ;
        RECT  0.33 0.33 2.20 59.75 ;
        RECT  0.33 108.90 2.20 109.60 ;
        RECT  0.33 241.90 2.20 242.60 ;
        RECT  0.33 380.90 2.20 559.92 ;
        RECT  14.70 0.33 103.70 559.92 ;

    END
END analog_gnd

MACRO analog_vdd
    CLASS PAD ;
    FOREIGN analog_vdd  0.00 -38.75 N  ;
    ORIGIN 0.00 39.15 ;
    SIZE 115.00 BY 600.00 ;
    SYMMETRY x y r90 ;
    SITE io_site ;
    PIN vdda!
        USE power ;  DIRECTION INOUT ;
        PORT
        CLASS CORE ;
        LAYER Metal1 ;
        RECT  14.00 -0.40 114.00 1.55 ;
        LAYER Metal2 ;
        RECT  14.00 -0.40 114.00 1.55 ;
        END
    END vdda!
    OBS
        LAYER Metal1 ;
        RECT  88.35 -0.40 114.75 560.00 ;
        RECT  86.55 0.90 88.35 560.00 ;
        RECT  0.25 -0.40 86.55 560.00 ;
        LAYER Metal2 ;
        RECT  0.33 0.33 114.68 559.92 ;
        LAYER Metal3 ;
        RECT  114.65 0.33 114.68 559.92 ;
        RECT  103.70 2.20 114.65 559.92 ;
        RECT  4.05 2.20 14.70 559.92 ;
        RECT  2.20 0.33 4.05 559.92 ;
        RECT  0.33 0.33 2.20 59.75 ;
        RECT  0.33 108.90 2.20 109.60 ;
        RECT  0.33 241.90 2.20 242.60 ;
        RECT  0.33 380.90 2.20 559.92 ;
        RECT  14.70 0.33 103.70 559.92 ;
        LAYER Metal4 ;
        RECT  0.33 0.33 114.68 559.92 ;
        LAYER Metal5 ;
        RECT  114.65 0.33 114.68 559.92 ;
        RECT  103.70 2.20 114.65 559.92 ;
        RECT  4.05 2.20 14.70 559.92 ;
        RECT  2.20 0.33 4.05 559.92 ;
        RECT  0.33 0.33 2.20 59.75 ;
        RECT  0.33 108.90 2.20 109.60 ;
        RECT  0.33 241.90 2.20 242.60 ;
        RECT  0.33 380.90 2.20 559.92 ;
        RECT  14.70 0.33 103.70 559.92 ;

    END
END analog_vdd



MACRO inbuf3_16pd
    CLASS PAD ;
    FOREIGN inbuf3_16pd  0.00 -38.75 N  ;
    ORIGIN 0.00 39.15 ;
    SIZE 115.00 BY 600.00 ;
    SYMMETRY x y r90 ;
    SITE io_site ;
    PIN di  USE SIGNAL ; DIRECTION OUTPUT ;
        PORT
        LAYER Metal1 ;
        RECT  87.15 -0.40 87.75 0.30 ;
        END
    END di
    PIN pad USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal3 ;
        RECT  3.00 383.00 112.00 544.25 ;
        END
    END pad
    PIN vdd!
        USE power ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        LAYER Metal3 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        END
    END vdd!
    PIN vss!
        USE ground ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        LAYER Metal3 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        END
    END vss!
    OBS
        LAYER Metal1 ;
        RECT  88.35 -0.40 114.75 560.00 ;
        RECT  86.55 0.90 88.35 560.00 ;
        RECT  0.25 -0.40 86.55 560.00 ;
        LAYER Metal2 ;
        RECT  0.33 0.33 114.68 559.92 ;
        LAYER Metal3 ;
        RECT  114.65 0.33 114.68 559.92 ;
        RECT  103.70 2.20 114.65 559.92 ;
        RECT  4.05 2.20 14.70 559.92 ;
        RECT  2.20 0.33 4.05 559.92 ;
        RECT  0.33 0.33 2.20 59.75 ;
        RECT  0.33 108.90 2.20 109.60 ;
        RECT  0.33 241.90 2.20 242.60 ;
        RECT  0.33 380.90 2.20 559.92 ;
        RECT  14.70 0.33 103.70 559.92 ;
    END
END inbuf3_16pd

MACRO inbuf3_16pu
    CLASS PAD ;
    FOREIGN inbuf3_16pu  0.00 -38.75 N  ;
    ORIGIN 0.00 39.15 ;
    SIZE 115.00 BY 600.00 ;
    SYMMETRY x y r90 ;
    SITE io_site ;
    PIN di  USE SIGNAL ; DIRECTION OUTPUT ;
        PORT
        LAYER Metal1 ;
        RECT  87.15 -0.40 87.75 0.30 ;
        END
    END di
    PIN pad USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal3 ;
        RECT  3.00 383.00 112.00 544.25 ;
        END
    END pad
    PIN vdd!
        USE power ;  DIRECTION INOUT ;
        PORT
        CLASS CORE ;
        LAYER Metal2 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        LAYER Metal3 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        END
    END vdd!
    PIN vss!
        USE ground ;  DIRECTION INOUT ;
        PORT
        CLASS CORE ;
        LAYER Metal2 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        LAYER Metal3 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        END
    END vss!
    OBS
        LAYER Metal1 ;
        RECT  88.35 -0.40 114.75 560.00 ;
        RECT  86.55 0.90 88.35 560.00 ;
        RECT  0.25 -0.40 86.55 560.00 ;
        LAYER Metal2 ;
        RECT  0.33 0.33 114.68 559.92 ;
        LAYER Metal3 ;
        RECT  114.65 0.33 114.68 559.92 ;
        RECT  103.70 2.20 114.65 559.92 ;
        RECT  4.05 2.20 14.70 559.92 ;
        RECT  2.20 0.33 4.05 559.92 ;
        RECT  0.33 0.33 2.20 59.75 ;
        RECT  0.33 108.90 2.20 109.60 ;
        RECT  0.33 241.90 2.20 242.60 ;
        RECT  0.33 380.90 2.20 559.92 ;
        RECT  14.70 0.33 103.70 559.92 ;
    END
END inbuf3_16pu

MACRO inbufs2_16
    CLASS PAD ;
    FOREIGN inbufs2_16  0.00 -38.75 N  ;
    ORIGIN 0.00 39.15 ;
    SIZE 115.00 BY 600.00 ;
    SYMMETRY x y r90 ;
    SITE io_site ;
    PIN di  USE SIGNAL ; DIRECTION OUTPUT ;
        PORT
        LAYER Metal1 ;
        RECT  87.15 -0.40 87.75 0.30 ;
        END
    END di
    PIN pad USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal3 ;
        RECT  3.00 383.00 112.00 544.25 ;
        END
    END pad
    PIN vdd!
        USE power ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        LAYER Metal3 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        END
    END vdd!
    PIN vss!
        USE ground ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        LAYER Metal3 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        END
    END vss!
    OBS
        LAYER Metal1 ;
        RECT  88.35 -0.40 114.75 560.00 ;
        RECT  86.55 0.90 88.35 560.00 ;
        RECT  0.25 -0.40 86.55 560.00 ;
        LAYER Metal2 ;
        RECT  0.33 0.33 114.68 559.92 ;
        LAYER Metal3 ;
        RECT  114.65 0.33 114.68 559.92 ;
        RECT  103.70 2.20 114.65 559.92 ;
        RECT  4.05 2.20 14.70 559.92 ;
        RECT  2.20 0.33 4.05 559.92 ;
        RECT  0.33 0.33 2.20 59.75 ;
        RECT  0.33 108.90 2.20 109.60 ;
        RECT  0.33 241.90 2.20 242.60 ;
        RECT  0.33 380.90 2.20 559.92 ;
        RECT  14.70 0.33 103.70 559.92 ;
    END
END inbufs2_16

MACRO inbufs2_16pd
    CLASS PAD ;
    FOREIGN inbufs2_16pd  0.00 -38.75 N  ;
    ORIGIN 0.00 39.15 ;
    SIZE 115.00 BY 600.00 ;
    SYMMETRY x y r90 ;
    SITE io_site ;
    PIN di  USE SIGNAL ; DIRECTION OUTPUT ;
        PORT
        LAYER Metal1 ;
        RECT  87.15 -0.40 87.75 0.30 ;
        END
    END di
    PIN pad USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal3 ;
        RECT  3.00 383.00 112.00 544.25 ;
        END
    END pad
    PIN vdd!
        USE power ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        LAYER Metal3 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        END
    END vdd!
    PIN vss!
        USE ground ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        LAYER Metal3 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        END
    END vss!
    OBS
        LAYER Metal1 ;
        RECT  88.35 -0.40 114.75 560.00 ;
        RECT  86.55 0.90 88.35 560.00 ;
        RECT  0.25 -0.40 86.55 560.00 ;
        LAYER Metal2 ;
        RECT  0.33 0.33 114.68 559.92 ;
        LAYER Metal3 ;
        RECT  114.65 0.33 114.68 559.92 ;
        RECT  103.70 2.20 114.65 559.92 ;
        RECT  4.05 2.20 14.70 559.92 ;
        RECT  2.20 0.33 4.05 559.92 ;
        RECT  0.33 0.33 2.20 59.75 ;
        RECT  0.33 108.90 2.20 109.60 ;
        RECT  0.33 241.90 2.20 242.60 ;
        RECT  0.33 380.90 2.20 559.92 ;
        RECT  14.70 0.33 103.70 559.92 ;
    END
END inbufs2_16pd

MACRO inbufs2_16pu
    CLASS PAD ;
    FOREIGN inbufs2_16pu  0.00 -38.75 N  ;
    ORIGIN 0.00 39.15 ;
    SIZE 115.00 BY 600.00 ;
    SYMMETRY x y r90 ;
    SITE io_site ;
    PIN di  USE SIGNAL ; DIRECTION OUTPUT ;
        PORT
        LAYER Metal1 ;
        RECT  87.15 -0.40 87.75 0.30 ;
        END
    END di
    PIN pad USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal3 ;
        RECT  3.00 383.00 112.00 544.25 ;
        END
    END pad
    PIN vdd!
        USE power ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        LAYER Metal3 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        END
    END vdd!
    PIN vss!
        USE ground ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        LAYER Metal3 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        END
    END vss!
    OBS
        LAYER Metal1 ;
        RECT  88.35 -0.40 114.75 560.00 ;
        RECT  86.55 0.90 88.35 560.00 ;
        RECT  0.25 -0.40 86.55 560.00 ;
        LAYER Metal2 ;
        RECT  0.33 0.33 114.68 559.92 ;
        LAYER Metal3 ;
        RECT  114.65 0.33 114.68 559.92 ;
        RECT  103.70 2.20 114.65 559.92 ;
        RECT  4.05 2.20 14.70 559.92 ;
        RECT  2.20 0.33 4.05 559.92 ;
        RECT  0.33 0.33 2.20 59.75 ;
        RECT  0.33 108.90 2.20 109.60 ;
        RECT  0.33 241.90 2.20 242.60 ;
        RECT  0.33 380.90 2.20 559.92 ;
        RECT  14.70 0.33 103.70 559.92 ;
    END
END inbufs2_16pu

MACRO inbufs3_16
    CLASS PAD ;
    FOREIGN inbufs3_16  0.00 -38.75 N  ;
    ORIGIN 0.00 39.15 ;
    SIZE 115.00 BY 600.00 ;
    SYMMETRY x y r90 ;
    SITE io_site ;
    PIN di  USE SIGNAL ; DIRECTION OUTPUT ;
        PORT
        LAYER Metal1 ;
        RECT  87.15 -0.40 87.75 0.30 ;
        END
    END di
    PIN pad USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal3 ;
        RECT  3.00 383.00 112.00 544.25 ;
        END
    END pad
    PIN vdd!
        USE power ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        LAYER Metal3 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        END
    END vdd!
    PIN vss!
        USE ground ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        LAYER Metal3 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        END
    END vss!
    OBS
        LAYER Metal1 ;
        RECT  88.35 -0.40 114.75 560.00 ;
        RECT  86.55 0.90 88.35 560.00 ;
        RECT  0.25 -0.40 86.55 560.00 ;
        LAYER Metal2 ;
        RECT  0.33 0.33 114.68 559.92 ;
        LAYER Metal3 ;
        RECT  114.65 0.33 114.68 559.92 ;
        RECT  103.70 2.20 114.65 559.92 ;
        RECT  4.05 2.20 14.70 559.92 ;
        RECT  2.20 0.33 4.05 559.92 ;
        RECT  0.33 0.33 2.20 59.75 ;
        RECT  0.33 108.90 2.20 109.60 ;
        RECT  0.33 241.90 2.20 242.60 ;
        RECT  0.33 380.90 2.20 559.92 ;
        RECT  14.70 0.33 103.70 559.92 ;
    END
END inbufs3_16

MACRO inbufs3_16pd
    CLASS PAD ;
    FOREIGN inbufs3_16pd  0.00 -38.75 N  ;
    ORIGIN 0.00 39.15 ;
    SIZE 115.00 BY 600.00 ;
    SYMMETRY x y r90 ;
    SITE io_site ;
    PIN di  USE SIGNAL ; DIRECTION OUTPUT ;
        PORT
        LAYER Metal1 ;
        RECT  87.15 -0.40 87.75 0.30 ;
        END
    END di
    PIN pad USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal3 ;
        RECT  3.00 383.00 112.00 544.25 ;
        END
    END pad
    PIN vdd!
        USE power ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        LAYER Metal3 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        END
    END vdd!
    PIN vss!
        USE ground ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        LAYER Metal3 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        END
    END vss!
    OBS
        LAYER Metal1 ;
        RECT  88.35 -0.40 114.75 560.00 ;
        RECT  86.55 0.90 88.35 560.00 ;
        RECT  0.25 -0.40 86.55 560.00 ;
        LAYER Metal2 ;
        RECT  0.33 0.33 114.68 559.92 ;
        LAYER Metal3 ;
        RECT  114.65 0.33 114.68 559.92 ;
        RECT  103.70 2.20 114.65 559.92 ;
        RECT  4.05 2.20 14.70 559.92 ;
        RECT  2.20 0.33 4.05 559.92 ;
        RECT  0.33 0.33 2.20 59.75 ;
        RECT  0.33 108.90 2.20 109.60 ;
        RECT  0.33 241.90 2.20 242.60 ;
        RECT  0.33 380.90 2.20 559.92 ;
        RECT  14.70 0.33 103.70 559.92 ;
    END
END inbufs3_16pd

MACRO inbufs3_16pu
    CLASS PAD ;
    FOREIGN inbufs3_16pu  0.00 -38.75 N  ;
    ORIGIN 0.00 39.15 ;
    SIZE 115.00 BY 600.00 ;
    SYMMETRY x y r90 ;
    SITE io_site ;
    PIN di  USE SIGNAL ; DIRECTION OUTPUT ;
        PORT
        LAYER Metal1 ;
        RECT  87.15 -0.40 87.75 0.30 ;
        END
    END di
    PIN pad USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal3 ;
        RECT  3.00 383.00 112.00 544.25 ;
        END
    END pad
    PIN vdd!
        USE power ;  DIRECTION INOUT ;
        PORT
        CLASS CORE ;
        LAYER Metal2 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        LAYER Metal3 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        END
    END vdd!
    PIN vss!
        USE ground ;  DIRECTION INOUT ;
        PORT
        CLASS CORE ;
        LAYER Metal2 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        LAYER Metal3 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        END
    END vss!
    OBS
        LAYER Metal1 ;
        RECT  88.35 -0.40 114.75 560.00 ;
        RECT  86.55 0.90 88.35 560.00 ;
        RECT  0.25 -0.40 86.55 560.00 ;
        LAYER Metal2 ;
        RECT  0.33 0.33 114.68 559.92 ;
        LAYER Metal3 ;
        RECT  114.65 0.33 114.68 559.92 ;
        RECT  103.70 2.20 114.65 559.92 ;
        RECT  4.05 2.20 14.70 559.92 ;
        RECT  2.20 0.33 4.05 559.92 ;
        RECT  0.33 0.33 2.20 59.75 ;
        RECT  0.33 108.90 2.20 109.60 ;
        RECT  0.33 241.90 2.20 242.60 ;
        RECT  0.33 380.90 2.20 559.92 ;
        RECT  14.70 0.33 103.70 559.92 ;
    END
END inbufs3_16pu

MACRO inpvdd
    CLASS PAD ;
    FOREIGN inpvdd  0.00 -38.75 N  ;
    ORIGIN 0.00 39.15 ;
    SIZE 115.00 BY 600.00 ;
    SYMMETRY x y r90 ;
    SITE io_site ;
    PIN pad USE POWER ; DIRECTION INPUT ;
        PORT
        LAYER Metal3 ;
        RECT  3.00 383.00 112.00 544.25 ;
        END
    END pad
    OBS
        LAYER Metal1 ;
        RECT  0.25 -0.40 114.75 560.00 ;
        LAYER Metal2 ;
        RECT  0.33 0.33 114.68 559.92 ;
        LAYER Metal3 ;
        RECT  0.33 0.33 114.68 559.92 ;
    END
END inpvdd

MACRO inpvss
    CLASS PAD ;
    FOREIGN inpvss  0.00 -38.75 N  ;
    ORIGIN 0.00 39.15 ;
    SIZE 115.00 BY 600.00 ;
    SYMMETRY x y r90 ;
    SITE io_site ;
    PIN pad USE power ; DIRECTION INPUT ;
        PORT
        LAYER Metal3 ;
        RECT  3.00 383.00 112.00 544.25 ;
        END
    END pad
    OBS
        LAYER Metal1 ;
        RECT  0.25 -0.40 114.75 560.00 ;
        LAYER Metal2 ;
        RECT  0.33 0.33 114.68 559.92 ;
        LAYER Metal3 ;
        RECT  0.33 0.33 114.68 559.92 ;
    END
END inpvss

MACRO io_fill_20
    CLASS PAD ;
    FOREIGN io_fill_20  0.00 -38.75 N  ;
    ORIGIN 0.00 39.15 ;
    SIZE 28.75 BY 600.00 ;
    SYMMETRY x y r90 ;
    SITE io_site ;
    OBS
        LAYER Metal1 ;
        RECT  0.25 -0.40 28.50 560.00 ;
        LAYER Metal2 ;
        RECT  0.33 0.33 28.43 559.92 ;
        LAYER Metal3 ;
        RECT  0.33 0.33 28.43 559.92 ;
        LAYER Metal4 ;
        RECT  0.33 0.33 28.43 559.92 ;
        LAYER Metal5 ;
        RECT  0.33 0.33 28.43 559.92 ;
    END
END io_fill_20

MACRO io_fill_40
    CLASS PAD ;
    FOREIGN io_fill_40  0.00 -38.75 N  ;
    ORIGIN 0.00 39.15 ;
    SIZE 57.50 BY 600.00 ;
    SYMMETRY x y r90 ;
    SITE io_site ;
    OBS
        LAYER Metal1 ;
        RECT  0.25 -0.40 57.16 560.00 ;
        LAYER Metal2 ;
        RECT  0.33 0.33 57.16 559.92 ;
        LAYER Metal3 ;
        RECT  0.33 0.33 57.16 559.92 ;
        LAYER Metal4 ;
        RECT  0.33 0.33 57.16 559.92 ;
        LAYER Metal5 ;
        RECT  0.33 0.33 57.16 559.92 ;
    END
END io_fill_40

MACRO io_fill_80
    CLASS PAD ;
    FOREIGN io_fill_80  0.00 -38.75 N  ;
    ORIGIN 0.00 39.15 ;
    SIZE 115.00 BY 600.00 ;
    SYMMETRY x y r90 ;
    SITE io_site ;
    OBS
        LAYER Metal1 ;
        RECT  0.25 -0.40 114.75 560.00 ;
        LAYER Metal2 ;
        RECT  0.33 0.33 114.67 559.92 ;
        LAYER Metal3 ;
        RECT  0.33 0.33 114.67 559.92 ;
        LAYER Metal4 ;
        RECT  0.33 0.33 114.67 559.92 ;
        LAYER Metal5 ;
        RECT  0.33 0.33 114.67 559.92 ;
    END
END io_fill_80

MACRO io_fill_80e
    CLASS PAD ;
    FOREIGN io_fill_80e  0.00 -38.75 N  ;
    ORIGIN 0.00 39.15 ;
    SIZE 115.00 BY 600.00 ;
    SYMMETRY x y r90 ;
    SITE io_site ;
    OBS
        LAYER Metal1 ;
        RECT  0.25 -0.40 114.75 560.00 ;
        LAYER Metal2 ;
        RECT  0.33 0.33 114.67 559.92 ;
        LAYER Metal3 ;
        RECT  0.33 0.33 114.67 559.92 ;
        LAYER Metal4 ;
        RECT  0.33 0.33 114.67 559.92 ;
        LAYER Metal5 ;
        RECT  0.33 0.33 114.67 559.92 ;
    END
END io_fill_80e

MACRO iobuf2_16_12
    CLASS PAD ;
    FOREIGN iobuf2_16_12  0.00 -38.75 N  ;
    ORIGIN 0.00 39.15 ;
    SIZE 115.00 BY 600.00 ;
    SYMMETRY x y r90 ;
    SITE io_site ;
     PIN en USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  60.95 -0.40 61.55 0.30 ;
        END
    END en
    PIN pad USE SIGNAL ; DIRECTION INOUT ;
        PORT
        LAYER Metal3 ;
        RECT  3.00 383.00 112.00 544.25 ;
        END
    END pad
    PIN do USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  25.95 -0.40 26.55 0.30 ;
        END
    END do
    PIN di  USE SIGNAL ; DIRECTION OUTPUT ;
        PORT
        LAYER Metal1 ;
        RECT  87.15 -0.40 87.75 0.30 ;
        END
    END di
    PIN vdd!
        USE power ;  DIRECTION INOUT ;
        PORT
        CLASS CORE ;
        LAYER Metal2 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        LAYER Metal3 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        END
    END vdd!
    PIN vss!
        USE ground ;  DIRECTION INOUT ;
        PORT
        CLASS CORE ;
        LAYER Metal2 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        LAYER Metal3 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        END
    END vss!
    OBS
        LAYER Metal1 ;
        RECT  88.35 -0.40 114.75 560.00 ;
        RECT  86.55 0.90 88.35 560.00 ;
        RECT  62.15 -0.40 86.55 560.00 ;
        RECT  60.35 0.90 62.15 560.00 ;
        RECT  27.15 -0.40 60.35 560.00 ;
        RECT  25.35 0.90 27.15 560.00 ;
        RECT  0.25 -0.40 25.35 560.00 ;
        LAYER Metal2 ;
        RECT  0.33 0.33 114.68 559.92 ;
        LAYER Metal3 ;
        RECT  114.65 0.33 114.68 559.92 ;
        RECT  103.70 2.20 114.65 559.92 ;
        RECT  4.05 2.20 14.70 559.92 ;
        RECT  2.20 0.33 4.05 559.92 ;
        RECT  0.33 0.33 2.20 59.75 ;
        RECT  0.33 108.90 2.20 109.60 ;
        RECT  0.33 241.90 2.20 242.60 ;
        RECT  0.33 380.90 2.20 559.92 ;
        RECT  14.70 0.33 103.70 559.92 ;
    END
END iobuf2_16_12

MACRO iobuf2_16_4
    CLASS PAD ;
    FOREIGN iobuf2_16_4  0.00 -38.75 N  ;
    ORIGIN 0.00 39.15 ;
    SIZE 115.00 BY 600.00 ;
    SYMMETRY x y r90 ;
    SITE io_site ;
     PIN en USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  60.95 -0.40 61.55 0.30 ;
        END
    END en
    PIN pad USE SIGNAL ; DIRECTION INOUT ;
        PORT
        LAYER Metal3 ;
        RECT  3.00 383.00 112.00 544.25 ;
        END
    END pad
    PIN do USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  25.95 -0.40 26.55 0.30 ;
        END
    END do
    PIN di  USE SIGNAL ; DIRECTION OUTPUT ;
        PORT
        LAYER Metal1 ;
        RECT  87.15 -0.40 87.75 0.30 ;
        END
    END di
    PIN vdd!
        USE power ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        LAYER Metal3 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        END
    END vdd!
    PIN vss!
        USE ground ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        LAYER Metal3 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        END
    END vss!
    OBS
        LAYER Metal1 ;
        RECT  88.35 -0.40 114.75 560.00 ;
        RECT  86.55 0.90 88.35 560.00 ;
        RECT  62.15 -0.40 86.55 560.00 ;
        RECT  60.35 0.90 62.15 560.00 ;
        RECT  27.15 -0.40 60.35 560.00 ;
        RECT  25.35 0.90 27.15 560.00 ;
        RECT  0.25 -0.40 25.35 560.00 ;
        LAYER Metal2 ;
        RECT  0.33 0.33 114.68 559.92 ;
        LAYER Metal3 ;
        RECT  114.65 0.33 114.68 559.92 ;
        RECT  103.70 2.20 114.65 559.92 ;
        RECT  4.05 2.20 14.70 559.92 ;
        RECT  2.20 0.33 4.05 559.92 ;
        RECT  0.33 0.33 2.20 59.75 ;
        RECT  0.33 108.90 2.20 109.60 ;
        RECT  0.33 241.90 2.20 242.60 ;
        RECT  0.33 380.90 2.20 559.92 ;
        RECT  14.70 0.33 103.70 559.92 ;
    END
END iobuf2_16_4

MACRO iobuf2_16_8
    CLASS PAD ;
    FOREIGN iobuf2_16_8  0.00 -38.75 N  ;
    ORIGIN 0.00 39.15 ;
    SIZE 115.00 BY 600.00 ;
    SYMMETRY x y r90 ;
    SITE io_site ;
     PIN en USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  60.95 -0.40 61.55 0.30 ;
        END
    END en
    PIN pad USE SIGNAL ; DIRECTION INOUT ;
        PORT
        LAYER Metal3 ;
        RECT  3.00 383.00 112.00 544.25 ;
        END
    END pad
    PIN do USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  25.95 -0.40 26.55 0.30 ;
        END
    END do
    PIN di  USE SIGNAL ; DIRECTION OUTPUT ;
        PORT
        LAYER Metal1 ;
        RECT  87.15 -0.40 87.75 0.30 ;
        END
    END di
    PIN vdd!
        USE power ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        LAYER Metal3 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        END
    END vdd!
    PIN vss!
        USE ground ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        LAYER Metal3 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        END
    END vss!
    OBS
        LAYER Metal1 ;
        RECT  88.35 -0.40 114.75 560.00 ;
        RECT  86.55 0.90 88.35 560.00 ;
        RECT  62.15 -0.40 86.55 560.00 ;
        RECT  60.35 0.90 62.15 560.00 ;
        RECT  27.15 -0.40 60.35 560.00 ;
        RECT  25.35 0.90 27.15 560.00 ;
        RECT  0.25 -0.40 25.35 560.00 ;
        LAYER Metal2 ;
        RECT  0.33 0.33 114.68 559.92 ;
        LAYER Metal3 ;
        RECT  114.65 0.33 114.68 559.92 ;
        RECT  103.70 2.20 114.65 559.92 ;
        RECT  4.05 2.20 14.70 559.92 ;
        RECT  2.20 0.33 4.05 559.92 ;
        RECT  0.33 0.33 2.20 59.75 ;
        RECT  0.33 108.90 2.20 109.60 ;
        RECT  0.33 241.90 2.20 242.60 ;
        RECT  0.33 380.90 2.20 559.92 ;
        RECT  14.70 0.33 103.70 559.92 ;
    END
END iobuf2_16_8

MACRO iobuf2_16pd_12
    CLASS PAD ;
    FOREIGN iobuf2_16pd_12  0.00 -38.75 N  ;
    ORIGIN 0.00 39.15 ;
    SIZE 115.00 BY 600.00 ;
    SYMMETRY x y r90 ;
    SITE io_site ;
     PIN en USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  60.95 -0.40 61.55 0.30 ;
        END
    END en
    PIN pad USE SIGNAL ; DIRECTION INOUT ;
        PORT
        LAYER Metal3 ;
        RECT  3.00 383.00 112.00 544.25 ;
        END
    END pad
    PIN do USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  25.95 -0.40 26.55 0.30 ;
        END
    END do
    PIN di  USE SIGNAL ; DIRECTION OUTPUT ;
        PORT
        LAYER Metal1 ;
        RECT  87.15 -0.40 87.75 0.30 ;
        END
    END di
    PIN vdd!
        USE power ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        LAYER Metal3 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        END
    END vdd!
    PIN vss!
        USE ground ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        LAYER Metal3 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        END
    END vss!
    OBS
        LAYER Metal1 ;
        RECT  88.35 -0.40 114.75 560.00 ;
        RECT  86.55 0.90 88.35 560.00 ;
        RECT  62.15 -0.40 86.55 560.00 ;
        RECT  60.35 0.90 62.15 560.00 ;
        RECT  27.15 -0.40 60.35 560.00 ;
        RECT  25.35 0.90 27.15 560.00 ;
        RECT  0.25 -0.40 25.35 560.00 ;
        LAYER Metal2 ;
        RECT  0.33 0.33 114.68 559.92 ;
        LAYER Metal3 ;
        RECT  114.65 0.33 114.68 559.92 ;
        RECT  103.70 2.20 114.65 559.92 ;
        RECT  4.05 2.20 14.70 559.92 ;
        RECT  2.20 0.33 4.05 559.92 ;
        RECT  0.33 0.33 2.20 59.75 ;
        RECT  0.33 108.90 2.20 109.60 ;
        RECT  0.33 241.90 2.20 242.60 ;
        RECT  0.33 380.90 2.20 559.92 ;
        RECT  14.70 0.33 103.70 559.92 ;
    END
END iobuf2_16pd_12

MACRO iobuf2_16pd_4
    CLASS PAD ;
    FOREIGN iobuf2_16pd_4  0.00 -38.75 N  ;
    ORIGIN 0.00 39.15 ;
    SIZE 115.00 BY 600.00 ;
    SYMMETRY x y r90 ;
    SITE io_site ;
     PIN en USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  60.95 -0.40 61.55 0.30 ;
        END
    END en
    PIN pad USE SIGNAL ; DIRECTION INOUT ;
        PORT
        LAYER Metal3 ;
        RECT  3.00 383.00 112.00 544.25 ;
        END
    END pad
    PIN do USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  25.95 -0.40 26.55 0.30 ;
        END
    END do
    PIN di  USE SIGNAL ; DIRECTION OUTPUT ;
        PORT
        LAYER Metal1 ;
        RECT  87.15 -0.40 87.75 0.30 ;
        END
    END di
    PIN vdd!
        USE power ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        LAYER Metal3 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        END
    END vdd!
    PIN vss!
        USE ground ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        LAYER Metal3 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        END
    END vss!
    OBS
        LAYER Metal1 ;
        RECT  88.35 -0.40 114.75 560.00 ;
        RECT  86.55 0.90 88.35 560.00 ;
        RECT  62.15 -0.40 86.55 560.00 ;
        RECT  60.35 0.90 62.15 560.00 ;
        RECT  27.15 -0.40 60.35 560.00 ;
        RECT  25.35 0.90 27.15 560.00 ;
        RECT  0.25 -0.40 25.35 560.00 ;
        LAYER Metal2 ;
        RECT  0.33 0.33 114.68 559.92 ;
        LAYER Metal3 ;
        RECT  114.65 0.33 114.68 559.92 ;
        RECT  103.70 2.20 114.65 559.92 ;
        RECT  4.05 2.20 14.70 559.92 ;
        RECT  2.20 0.33 4.05 559.92 ;
        RECT  0.33 0.33 2.20 59.75 ;
        RECT  0.33 108.90 2.20 109.60 ;
        RECT  0.33 241.90 2.20 242.60 ;
        RECT  0.33 380.90 2.20 559.92 ;
        RECT  14.70 0.33 103.70 559.92 ;
    END
END iobuf2_16pd_4

MACRO iobuf2_16pd_8
    CLASS PAD ;
    FOREIGN iobuf2_16pd_8  0.00 -38.75 N  ;
    ORIGIN 0.00 39.15 ;
    SIZE 115.00 BY 600.00 ;
    SYMMETRY x y r90 ;
    SITE io_site ;
     PIN en USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  60.95 -0.40 61.55 0.30 ;
        END
    END en
    PIN pad USE SIGNAL ; DIRECTION INOUT ;
        PORT
        LAYER Metal3 ;
        RECT  3.00 383.00 112.00 544.25 ;
        END
    END pad
    PIN do USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  25.95 -0.40 26.55 0.30 ;
        END
    END do
    PIN di  USE SIGNAL ; DIRECTION OUTPUT ;
        PORT
        LAYER Metal1 ;
        RECT  87.15 -0.40 87.75 0.30 ;
        END
    END di
    PIN vdd!
        USE power ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        LAYER Metal3 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        END
    END vdd!
    PIN vss!
        USE ground ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        LAYER Metal3 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        END
    END vss!
    OBS
        LAYER Metal1 ;
        RECT  88.35 -0.40 114.75 560.00 ;
        RECT  86.55 0.90 88.35 560.00 ;
        RECT  62.15 -0.40 86.55 560.00 ;
        RECT  60.35 0.90 62.15 560.00 ;
        RECT  27.15 -0.40 60.35 560.00 ;
        RECT  25.35 0.90 27.15 560.00 ;
        RECT  0.25 -0.40 25.35 560.00 ;
        LAYER Metal2 ;
        RECT  0.33 0.33 114.68 559.92 ;
        LAYER Metal3 ;
        RECT  114.65 0.33 114.68 559.92 ;
        RECT  103.70 2.20 114.65 559.92 ;
        RECT  4.05 2.20 14.70 559.92 ;
        RECT  2.20 0.33 4.05 559.92 ;
        RECT  0.33 0.33 2.20 59.75 ;
        RECT  0.33 108.90 2.20 109.60 ;
        RECT  0.33 241.90 2.20 242.60 ;
        RECT  0.33 380.90 2.20 559.92 ;
        RECT  14.70 0.33 103.70 559.92 ;
    END
END iobuf2_16pd_8

MACRO iobuf2_16pu_12
    CLASS PAD ;
    FOREIGN iobuf2_16pu_12  0.00 -38.75 N  ;
    ORIGIN 0.00 39.15 ;
    SIZE 115.00 BY 600.00 ;
    SYMMETRY x y r90 ;
    SITE io_site ;
     PIN en USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  60.95 -0.40 61.55 0.30 ;
        END
    END en
    PIN pad USE SIGNAL ; DIRECTION INOUT ;
        PORT
        LAYER Metal3 ;
        RECT  3.00 383.00 112.00 544.25 ;
        END
    END pad
    PIN do USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  25.95 -0.40 26.55 0.30 ;
        END
    END do
    PIN di  USE SIGNAL ; DIRECTION OUTPUT ;
        PORT
        LAYER Metal1 ;
        RECT  87.15 -0.40 87.75 0.30 ;
        END
    END di
    PIN vdd!
        USE power ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        LAYER Metal3 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        END
    END vdd!
    PIN vss!
        USE ground ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        LAYER Metal3 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        END
    END vss!
    OBS
        LAYER Metal1 ;
        RECT  88.35 -0.40 114.75 560.00 ;
        RECT  86.55 0.90 88.35 560.00 ;
        RECT  62.15 -0.40 86.55 560.00 ;
        RECT  60.35 0.90 62.15 560.00 ;
        RECT  27.15 -0.40 60.35 560.00 ;
        RECT  25.35 0.90 27.15 560.00 ;
        RECT  0.25 -0.40 25.35 560.00 ;
        LAYER Metal2 ;
        RECT  0.33 0.33 114.68 559.92 ;
        LAYER Metal3 ;
        RECT  114.65 0.33 114.68 559.92 ;
        RECT  103.70 2.20 114.65 559.92 ;
        RECT  4.05 2.20 14.70 559.92 ;
        RECT  2.20 0.33 4.05 559.92 ;
        RECT  0.33 0.33 2.20 59.75 ;
        RECT  0.33 108.90 2.20 109.60 ;
        RECT  0.33 241.90 2.20 242.60 ;
        RECT  0.33 380.90 2.20 559.92 ;
        RECT  14.70 0.33 103.70 559.92 ;
    END
END iobuf2_16pu_12

MACRO iobuf2_16pu_4
    CLASS PAD ;
    FOREIGN iobuf2_16pu_4  0.00 -38.75 N  ;
    ORIGIN 0.00 39.15 ;
    SIZE 115.00 BY 600.00 ;
    SYMMETRY x y r90 ;
    SITE io_site ;
     PIN en USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  60.95 -0.40 61.55 0.30 ;
        END
    END en
    PIN pad USE SIGNAL ; DIRECTION INOUT ;
        PORT
        LAYER Metal3 ;
        RECT  3.00 383.00 112.00 544.25 ;
        END
    END pad
    PIN do USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  25.95 -0.40 26.55 0.30 ;
        END
    END do
    PIN di  USE SIGNAL ; DIRECTION OUTPUT ;
        PORT
        LAYER Metal1 ;
        RECT  87.15 -0.40 87.75 0.30 ;
        END
    END di
    PIN vdd!
        USE power ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        LAYER Metal3 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        END
    END vdd!
    PIN vss!
        USE ground ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        LAYER Metal3 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        END
    END vss!
    OBS
        LAYER Metal1 ;
        RECT  88.35 -0.40 114.75 560.00 ;
        RECT  86.55 0.90 88.35 560.00 ;
        RECT  62.15 -0.40 86.55 560.00 ;
        RECT  60.35 0.90 62.15 560.00 ;
        RECT  27.15 -0.40 60.35 560.00 ;
        RECT  25.35 0.90 27.15 560.00 ;
        RECT  0.25 -0.40 25.35 560.00 ;
        LAYER Metal2 ;
        RECT  0.33 0.33 114.68 559.92 ;
        LAYER Metal3 ;
        RECT  114.65 0.33 114.68 559.92 ;
        RECT  103.70 2.20 114.65 559.92 ;
        RECT  4.05 2.20 14.70 559.92 ;
        RECT  2.20 0.33 4.05 559.92 ;
        RECT  0.33 0.33 2.20 59.75 ;
        RECT  0.33 108.90 2.20 109.60 ;
        RECT  0.33 241.90 2.20 242.60 ;
        RECT  0.33 380.90 2.20 559.92 ;
        RECT  14.70 0.33 103.70 559.92 ;
    END
END iobuf2_16pu_4

MACRO iobuf2_16pu_8
    CLASS PAD ;
    FOREIGN iobuf2_16pu_8  0.00 -38.75 N  ;
    ORIGIN 0.00 39.15 ;
    SIZE 115.00 BY 600.00 ;
    SYMMETRY x y r90 ;
    SITE io_site ;
     PIN en USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  60.95 -0.40 61.55 0.30 ;
        END
    END en
    PIN pad USE SIGNAL ; DIRECTION INOUT ;
        PORT
        LAYER Metal3 ;
        RECT  3.00 383.00 112.00 544.25 ;
        END
    END pad
    PIN do USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  25.95 -0.40 26.55 0.30 ;
        END
    END do
    PIN di  USE SIGNAL ; DIRECTION OUTPUT ;
        PORT
        LAYER Metal1 ;
        RECT  87.15 -0.40 87.75 0.30 ;
        END
    END di
    PIN vdd!
        USE power ;  DIRECTION INOUT ;
        PORT
        CLASS CORE ;
        LAYER Metal2 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        LAYER Metal3 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        END
    END vdd!
    PIN vss!
        USE ground ;  DIRECTION INOUT ;
        PORT
        CLASS CORE ;
        LAYER Metal2 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        LAYER Metal3 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        END
    END vss!
    OBS
        LAYER Metal1 ;
        RECT  88.35 -0.40 114.75 560.00 ;
        RECT  86.55 0.90 88.35 560.00 ;
        RECT  62.15 -0.40 86.55 560.00 ;
        RECT  60.35 0.90 62.15 560.00 ;
        RECT  27.15 -0.40 60.35 560.00 ;
        RECT  25.35 0.90 27.15 560.00 ;
        RECT  0.25 -0.40 25.35 560.00 ;
        LAYER Metal2 ;
        RECT  0.33 0.33 114.68 559.92 ;
        LAYER Metal3 ;
        RECT  114.65 0.33 114.68 559.92 ;
        RECT  103.70 2.20 114.65 559.92 ;
        RECT  4.05 2.20 14.70 559.92 ;
        RECT  2.20 0.33 4.05 559.92 ;
        RECT  0.33 0.33 2.20 59.75 ;
        RECT  0.33 108.90 2.20 109.60 ;
        RECT  0.33 241.90 2.20 242.60 ;
        RECT  0.33 380.90 2.20 559.92 ;
        RECT  14.70 0.33 103.70 559.92 ;
    END
END iobuf2_16pu_8

MACRO iobuf3_16_12
    CLASS PAD ;
    FOREIGN iobuf3_16_12  0.00 -38.75 N  ;
    ORIGIN 0.00 39.15 ;
    SIZE 115.00 BY 600.00 ;
    SYMMETRY x y r90 ;
    SITE io_site ;
     PIN en USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  60.95 -0.40 61.55 0.30 ;
        END
    END en
    PIN pad USE SIGNAL ; DIRECTION INOUT ;
        PORT
        LAYER Metal5 ;
        RECT  3.00 383.00 112.00 544.25 ;
        END
    END pad
    PIN do USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  25.95 -0.40 26.55 0.30 ;
        END
    END do
    PIN di  USE SIGNAL ; DIRECTION OUTPUT ;
        PORT
        LAYER Metal1 ;
        RECT  87.15 -0.40 87.75 0.30 ;
        END
    END di
    PIN vdd!
        USE power ;  DIRECTION INOUT ;
        PORT
        CLASS CORE ;
        LAYER Metal2 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        LAYER Metal3 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        END
    END vdd!
    PIN vss!
        USE ground ;  DIRECTION INOUT ;
        PORT
        CLASS CORE ;
        LAYER Metal2 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        LAYER Metal3 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        END
    END vss!
    OBS
        LAYER Metal1 ;
        RECT  88.35 -0.40 114.75 560.00 ;
        RECT  86.55 0.90 88.35 560.00 ;
        RECT  62.15 -0.40 86.55 560.00 ;
        RECT  60.35 0.90 62.15 560.00 ;
        RECT  27.15 -0.40 60.35 560.00 ;
        RECT  25.35 0.90 27.15 560.00 ;
        RECT  0.25 -0.40 25.35 560.00 ;
        LAYER Metal2 ;
        RECT  0.33 0.33 114.68 559.92 ;
        LAYER Metal3 ;
        RECT  114.65 0.33 114.68 559.92 ;
        RECT  103.70 2.20 114.65 559.92 ;
        RECT  4.05 2.20 14.70 559.92 ;
        RECT  2.20 0.33 4.05 559.92 ;
        RECT  0.33 0.33 2.20 59.75 ;
        RECT  0.33 108.90 2.20 109.60 ;
        RECT  0.33 241.90 2.20 242.60 ;
        RECT  0.33 380.90 2.20 559.92 ;
        RECT  14.70 0.33 103.70 559.92 ;
        LAYER Metal4 ;
        RECT  0.33 0.33 114.68 559.92 ;
        LAYER Metal5 ;
        RECT  114.65 0.33 114.68 559.92 ;
        RECT  103.70 2.20 114.65 559.92 ;
        RECT  4.05 2.20 14.70 559.92 ;
        RECT  2.20 0.33 4.05 559.92 ;
        RECT  0.33 0.33 2.20 59.75 ;
        RECT  0.33 108.90 2.20 109.60 ;
        RECT  0.33 241.90 2.20 242.60 ;
        RECT  0.33 380.90 2.20 559.92 ;
        RECT  14.70 0.33 103.70 559.92 ;
    END
END iobuf3_16_12

MACRO iobuf3_16_4
    CLASS PAD ;
    FOREIGN iobuf3_16_4  0.00 -38.75 N  ;
    ORIGIN 0.00 39.15 ;
    SIZE 115.00 BY 600.00 ;
    SYMMETRY x y r90 ;
    SITE io_site ;
     PIN en USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  60.95 -0.40 61.55 0.30 ;
        END
    END en
    PIN pad USE SIGNAL ; DIRECTION INOUT ;
        PORT
        LAYER Metal3 ;
        RECT  3.00 383.00 112.00 544.25 ;
        END
    END pad
    PIN do USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  25.95 -0.40 26.55 0.30 ;
        END
    END do
    PIN di  USE SIGNAL ; DIRECTION OUTPUT ;
        PORT
        LAYER Metal1 ;
        RECT  87.15 -0.40 87.75 0.30 ;
        END
    END di
    PIN vdd!
        USE power ;  DIRECTION INOUT ;
        PORT
        CLASS CORE ;
        LAYER Metal2 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        LAYER Metal3 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        END
    END vdd!
    PIN vss!
        USE ground ;  DIRECTION INOUT ;
        PORT
        CLASS CORE ;
        LAYER Metal2 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        LAYER Metal3 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        END
    END vss!
    OBS
        LAYER Metal1 ;
        RECT  88.35 -0.40 114.75 560.00 ;
        RECT  86.55 0.90 88.35 560.00 ;
        RECT  62.15 -0.40 86.55 560.00 ;
        RECT  60.35 0.90 62.15 560.00 ;
        RECT  27.15 -0.40 60.35 560.00 ;
        RECT  25.35 0.90 27.15 560.00 ;
        RECT  0.25 -0.40 25.35 560.00 ;
        LAYER Metal2 ;
        RECT  0.33 0.33 114.68 559.92 ;
        LAYER Metal3 ;
        RECT  114.65 0.33 114.68 559.92 ;
        RECT  103.70 2.20 114.65 559.92 ;
        RECT  4.05 2.20 14.70 559.92 ;
        RECT  2.20 0.33 4.05 559.92 ;
        RECT  0.33 0.33 2.20 59.75 ;
        RECT  0.33 108.90 2.20 109.60 ;
        RECT  0.33 241.90 2.20 242.60 ;
        RECT  0.33 380.90 2.20 559.92 ;
        RECT  14.70 0.33 103.70 559.92 ;
    END
END iobuf3_16_4

MACRO iobuf3_16_8
    CLASS PAD ;
    FOREIGN iobuf3_16_8  0.00 -38.75 N  ;
    ORIGIN 0.00 39.15 ;
    SIZE 115.00 BY 600.00 ;
    SYMMETRY x y r90 ;
    SITE io_site ;
     PIN en USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  60.95 -0.40 61.55 0.30 ;
        END
    END en
    PIN pad USE SIGNAL ; DIRECTION INOUT ;
        PORT
        LAYER Metal5 ;
        RECT  3.00 383.00 112.00 544.25 ;
        END
    END pad
    PIN do USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  25.95 -0.40 26.55 0.30 ;
        END
    END do
    PIN di  USE SIGNAL ; DIRECTION OUTPUT ;
        PORT
        LAYER Metal1 ;
        RECT  87.15 -0.40 87.75 0.30 ;
        END
    END di
    PIN vdd!
        USE power ;  DIRECTION INOUT ;
        PORT
        CLASS CORE ;
        LAYER Metal2 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        LAYER Metal3 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        END
    END vdd!
    PIN vss!
        USE ground ;  DIRECTION INOUT ;
        PORT
        CLASS CORE ;
        LAYER Metal2 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        LAYER Metal3 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        END
    END vss!
    OBS
        LAYER Metal1 ;
        RECT  88.35 -0.40 114.75 560.00 ;
        RECT  86.55 0.90 88.35 560.00 ;
        RECT  62.15 -0.40 86.55 560.00 ;
        RECT  60.35 0.90 62.15 560.00 ;
        RECT  27.15 -0.40 60.35 560.00 ;
        RECT  25.35 0.90 27.15 560.00 ;
        RECT  0.25 -0.40 25.35 560.00 ;
        LAYER Metal2 ;
        RECT  0.33 0.33 114.68 559.92 ;
        LAYER Metal3 ;
        RECT  114.65 0.33 114.68 559.92 ;
        RECT  103.70 2.20 114.65 559.92 ;
        RECT  4.05 2.20 14.70 559.92 ;
        RECT  2.20 0.33 4.05 559.92 ;
        RECT  0.33 0.33 2.20 59.75 ;
        RECT  0.33 108.90 2.20 109.60 ;
        RECT  0.33 241.90 2.20 242.60 ;
        RECT  0.33 380.90 2.20 559.92 ;
        RECT  14.70 0.33 103.70 559.92 ;
        LAYER Metal4 ;
        RECT  0.33 0.33 114.68 559.92 ;
        LAYER Metal5 ;
        RECT  114.65 0.33 114.68 559.92 ;
        RECT  103.70 2.20 114.65 559.92 ;
        RECT  4.05 2.20 14.70 559.92 ;
        RECT  2.20 0.33 4.05 559.92 ;
        RECT  0.33 0.33 2.20 59.75 ;
        RECT  0.33 108.90 2.20 109.60 ;
        RECT  0.33 241.90 2.20 242.60 ;
        RECT  0.33 380.90 2.20 559.92 ;
        RECT  14.70 0.33 103.70 559.92 ;

    END
END iobuf3_16_8

MACRO iobuf3_16pd_12
    CLASS PAD ;
    FOREIGN iobuf3_16pd_12  0.00 -38.75 N  ;
    ORIGIN 0.00 39.15 ;
    SIZE 115.00 BY 600.00 ;
    SYMMETRY x y r90 ;
    SITE io_site ;
     PIN en USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  60.95 -0.40 61.55 0.30 ;
        END
    END en
    PIN pad USE SIGNAL ; DIRECTION INOUT ;
        PORT
        LAYER Metal3 ;
        RECT  3.00 383.00 112.00 544.25 ;
        END
    END pad
    PIN do USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  25.95 -0.40 26.55 0.30 ;
        END
    END do
    PIN di  USE SIGNAL ; DIRECTION OUTPUT ;
        PORT
        LAYER Metal1 ;
        RECT  87.15 -0.40 87.75 0.30 ;
        END
    END di
    PIN vdd!
        USE power ;  DIRECTION INOUT ;
        PORT
        CLASS CORE ;
        LAYER Metal2 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        LAYER Metal3 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        END
    END vdd!
    PIN vss!
        USE ground ;  DIRECTION INOUT ;
        PORT
        CLASS CORE ;
        LAYER Metal2 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        LAYER Metal3 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        END
    END vss!
    OBS
        LAYER Metal1 ;
        RECT  88.35 -0.40 114.75 560.00 ;
        RECT  86.55 0.90 88.35 560.00 ;
        RECT  62.15 -0.40 86.55 560.00 ;
        RECT  60.35 0.90 62.15 560.00 ;
        RECT  27.15 -0.40 60.35 560.00 ;
        RECT  25.35 0.90 27.15 560.00 ;
        RECT  0.25 -0.40 25.35 560.00 ;
        LAYER Metal2 ;
        RECT  0.33 0.33 114.68 559.92 ;
        LAYER Metal3 ;
        RECT  114.65 0.33 114.68 559.92 ;
        RECT  103.70 2.20 114.65 559.92 ;
        RECT  4.05 2.20 14.70 559.92 ;
        RECT  2.20 0.33 4.05 559.92 ;
        RECT  0.33 0.33 2.20 59.75 ;
        RECT  0.33 108.90 2.20 109.60 ;
        RECT  0.33 241.90 2.20 242.60 ;
        RECT  0.33 380.90 2.20 559.92 ;
        RECT  14.70 0.33 103.70 559.92 ;
    END
END iobuf3_16pd_12

MACRO iobuf3_16pd_4
    CLASS PAD ;
    FOREIGN iobuf3_16pd_4  0.00 -38.75 N  ;
    ORIGIN 0.00 39.15 ;
    SIZE 115.00 BY 600.00 ;
    SYMMETRY x y r90 ;
    SITE io_site ;
     PIN en USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  60.95 -0.40 61.55 0.30 ;
        END
    END en
    PIN pad USE SIGNAL ; DIRECTION INOUT ;
        PORT
        LAYER Metal3 ;
        RECT  3.00 383.00 112.00 544.25 ;
        END
    END pad
    PIN do USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  25.95 -0.40 26.55 0.30 ;
        END
    END do
    PIN di  USE SIGNAL ; DIRECTION OUTPUT ;
        PORT
        LAYER Metal1 ;
        RECT  87.15 -0.40 87.75 0.30 ;
        END
    END di
    PIN vdd!
        USE power ;  DIRECTION INOUT ;
        PORT
        CLASS CORE ;
        LAYER Metal2 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        LAYER Metal3 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        END
    END vdd!
    PIN vss!
        USE ground ;  DIRECTION INOUT ;
        PORT
        CLASS CORE ;
        LAYER Metal2 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        LAYER Metal3 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        END
    END vss!
    OBS
        LAYER Metal1 ;
        RECT  88.35 -0.40 114.75 560.00 ;
        RECT  86.55 0.90 88.35 560.00 ;
        RECT  62.15 -0.40 86.55 560.00 ;
        RECT  60.35 0.90 62.15 560.00 ;
        RECT  27.15 -0.40 60.35 560.00 ;
        RECT  25.35 0.90 27.15 560.00 ;
        RECT  0.25 -0.40 25.35 560.00 ;
        LAYER Metal2 ;
        RECT  0.33 0.33 114.68 559.92 ;
        LAYER Metal3 ;
        RECT  114.65 0.33 114.68 559.92 ;
        RECT  103.70 2.20 114.65 559.92 ;
        RECT  4.05 2.20 14.70 559.92 ;
        RECT  2.20 0.33 4.05 559.92 ;
        RECT  0.33 0.33 2.20 59.75 ;
        RECT  0.33 108.90 2.20 109.60 ;
        RECT  0.33 241.90 2.20 242.60 ;
        RECT  0.33 380.90 2.20 559.92 ;
        RECT  14.70 0.33 103.70 559.92 ;
    END
END iobuf3_16pd_4

MACRO iobuf3_16pd_8
    CLASS PAD ;
    FOREIGN iobuf3_16pd_8  0.00 -38.75 N  ;
    ORIGIN 0.00 39.15 ;
    SIZE 115.00 BY 600.00 ;
    SYMMETRY x y r90 ;
    SITE io_site ;
     PIN en USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  60.95 -0.40 61.55 0.30 ;
        END
    END en
    PIN pad USE SIGNAL ; DIRECTION INOUT ;
        PORT
        LAYER Metal3 ;
        RECT  3.00 383.00 112.00 544.25 ;
        END
    END pad
    PIN do USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  25.95 -0.40 26.55 0.30 ;
        END
    END do
    PIN di  USE SIGNAL ; DIRECTION OUTPUT ;
        PORT
        LAYER Metal1 ;
        RECT  87.15 -0.40 87.75 0.30 ;
        END
    END di
    PIN vdd!
        USE power ;  DIRECTION INOUT ;
        PORT
        CLASS CORE ;
        LAYER Metal2 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        LAYER Metal3 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        END
    END vdd!
    PIN vss!
        USE ground ;  DIRECTION INOUT ;
        PORT
        CLASS CORE ;
        LAYER Metal2 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        LAYER Metal3 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        END
    END vss!
    OBS
        LAYER Metal1 ;
        RECT  88.35 -0.40 114.75 560.00 ;
        RECT  86.55 0.90 88.35 560.00 ;
        RECT  62.15 -0.40 86.55 560.00 ;
        RECT  60.35 0.90 62.15 560.00 ;
        RECT  27.15 -0.40 60.35 560.00 ;
        RECT  25.35 0.90 27.15 560.00 ;
        RECT  0.25 -0.40 25.35 560.00 ;
        LAYER Metal2 ;
        RECT  0.33 0.33 114.68 559.92 ;
        LAYER Metal3 ;
        RECT  114.65 0.33 114.68 559.92 ;
        RECT  103.70 2.20 114.65 559.92 ;
        RECT  4.05 2.20 14.70 559.92 ;
        RECT  2.20 0.33 4.05 559.92 ;
        RECT  0.33 0.33 2.20 59.75 ;
        RECT  0.33 108.90 2.20 109.60 ;
        RECT  0.33 241.90 2.20 242.60 ;
        RECT  0.33 380.90 2.20 559.92 ;
        RECT  14.70 0.33 103.70 559.92 ;
    END
END iobuf3_16pd_8

MACRO iobuf3_16pu_12
    CLASS PAD ;
    FOREIGN iobuf3_16pu_12  0.00 -38.75 N  ;
    ORIGIN 0.00 39.15 ;
    SIZE 115.00 BY 600.00 ;
    SYMMETRY x y r90 ;
    SITE io_site ;
     PIN en USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  60.95 -0.40 61.55 0.30 ;
        END
    END en
    PIN pad USE SIGNAL ; DIRECTION INOUT ;
        PORT
        LAYER Metal3 ;
        RECT  3.00 383.00 112.00 544.25 ;
        END
    END pad
    PIN do USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  25.95 -0.40 26.55 0.30 ;
        END
    END do
    PIN di  USE SIGNAL ; DIRECTION OUTPUT ;
        PORT
        LAYER Metal1 ;
        RECT  87.15 -0.40 87.75 0.30 ;
        END
    END di
    PIN vdd!
        USE power ;  DIRECTION INOUT ;
        PORT
        CLASS CORE ;
        LAYER Metal2 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        LAYER Metal3 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        END
    END vdd!
    PIN vss!
        USE ground ;  DIRECTION INOUT ;
        PORT
        CLASS CORE ;
        LAYER Metal2 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        LAYER Metal3 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        END
    END vss!
    OBS
        LAYER Metal1 ;
        RECT  88.35 -0.40 114.75 560.00 ;
        RECT  86.55 0.90 88.35 560.00 ;
        RECT  62.15 -0.40 86.55 560.00 ;
        RECT  60.35 0.90 62.15 560.00 ;
        RECT  27.15 -0.40 60.35 560.00 ;
        RECT  25.35 0.90 27.15 560.00 ;
        RECT  0.25 -0.40 25.35 560.00 ;
        LAYER Metal2 ;
        RECT  0.33 0.33 114.68 559.92 ;
        LAYER Metal3 ;
        RECT  114.65 0.33 114.68 559.92 ;
        RECT  103.70 2.20 114.65 559.92 ;
        RECT  4.05 2.20 14.70 559.92 ;
        RECT  2.20 0.33 4.05 559.92 ;
        RECT  0.33 0.33 2.20 59.75 ;
        RECT  0.33 108.90 2.20 109.60 ;
        RECT  0.33 241.90 2.20 242.60 ;
        RECT  0.33 380.90 2.20 559.92 ;
        RECT  14.70 0.33 103.70 559.92 ;
    END
END iobuf3_16pu_12

MACRO iobuf3_16pu_4
    CLASS PAD ;
    FOREIGN iobuf3_16pu_4  0.00 -38.75 N  ;
    ORIGIN 0.00 39.15 ;
    SIZE 115.00 BY 600.00 ;
    SYMMETRY x y r90 ;
    SITE io_site ;
     PIN en USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  60.95 -0.40 61.55 0.30 ;
        END
    END en
    PIN pad USE SIGNAL ; DIRECTION INOUT ;
        PORT
        LAYER Metal3 ;
        RECT  3.00 383.00 112.00 544.25 ;
        END
    END pad
    PIN do USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  25.95 -0.40 26.55 0.30 ;
        END
    END do
    PIN di  USE SIGNAL ; DIRECTION OUTPUT ;
        PORT
        LAYER Metal1 ;
        RECT  87.15 -0.40 87.75 0.30 ;
        END
    END di
    PIN vdd!
        USE power ;  DIRECTION INOUT ;
        PORT
        CLASS CORE ;
        LAYER Metal2 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        LAYER Metal3 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        END
    END vdd!
    PIN vss!
        USE ground ;  DIRECTION INOUT ;
        PORT
        CLASS CORE ;
        LAYER Metal2 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        LAYER Metal3 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        END
    END vss!
    OBS
        LAYER Metal1 ;
        RECT  88.35 -0.40 114.75 560.00 ;
        RECT  86.55 0.90 88.35 560.00 ;
        RECT  62.15 -0.40 86.55 560.00 ;
        RECT  60.35 0.90 62.15 560.00 ;
        RECT  27.15 -0.40 60.35 560.00 ;
        RECT  25.35 0.90 27.15 560.00 ;
        RECT  0.25 -0.40 25.35 560.00 ;
        LAYER Metal2 ;
        RECT  0.33 0.33 114.68 559.92 ;
        LAYER Metal3 ;
        RECT  114.65 0.33 114.68 559.92 ;
        RECT  103.70 2.20 114.65 559.92 ;
        RECT  4.05 2.20 14.70 559.92 ;
        RECT  2.20 0.33 4.05 559.92 ;
        RECT  0.33 0.33 2.20 59.75 ;
        RECT  0.33 108.90 2.20 109.60 ;
        RECT  0.33 241.90 2.20 242.60 ;
        RECT  0.33 380.90 2.20 559.92 ;
        RECT  14.70 0.33 103.70 559.92 ;
    END
END iobuf3_16pu_4

MACRO iobuf3_16pu_8
    CLASS PAD ;
    FOREIGN iobuf3_16pu_8  0.00 -38.75 N  ;
    ORIGIN 0.00 39.15 ;
    SIZE 115.00 BY 600.00 ;
    SYMMETRY x y r90 ;
    SITE io_site ;
     PIN en USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  60.95 -0.40 61.55 0.30 ;
        END
    END en
    PIN pad USE SIGNAL ; DIRECTION INOUT ;
        PORT
        LAYER Metal5 ;
        RECT  3.00 383.00 112.00 544.25 ;
        END
    END pad
    PIN do USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  25.95 -0.40 26.55 0.30 ;
        END
    END do
    PIN di  USE SIGNAL ; DIRECTION OUTPUT ;
        PORT
        LAYER Metal1 ;
        RECT  87.15 -0.40 87.75 0.30 ;
        END
    END di
    PIN vdd!
        USE power ;  DIRECTION INOUT ;
        PORT
        CLASS CORE ;
        LAYER Metal2 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        LAYER Metal3 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        END
    END vdd!
    PIN vss!
        USE ground ;  DIRECTION INOUT ;
        PORT
        CLASS CORE ;
        LAYER Metal2 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        LAYER Metal3 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        END
    END vss!
    OBS
        LAYER Metal1 ;
        RECT  88.35 -0.40 114.75 560.00 ;
        RECT  86.55 0.90 88.35 560.00 ;
        RECT  62.15 -0.40 86.55 560.00 ;
        RECT  60.35 0.90 62.15 560.00 ;
        RECT  27.15 -0.40 60.35 560.00 ;
        RECT  25.35 0.90 27.15 560.00 ;
        RECT  0.25 -0.40 25.35 560.00 ;
        LAYER Metal2 ;
        RECT  0.33 0.33 114.68 559.92 ;
        LAYER Metal3 ;
        RECT  114.65 0.33 114.68 559.92 ;
        RECT  103.70 2.20 114.65 559.92 ;
        RECT  4.05 2.20 14.70 559.92 ;
        RECT  2.20 0.33 4.05 559.92 ;
        RECT  0.33 0.33 2.20 59.75 ;
        RECT  0.33 108.90 2.20 109.60 ;
        RECT  0.33 241.90 2.20 242.60 ;
        RECT  0.33 380.90 2.20 559.92 ;
        RECT  14.70 0.33 103.70 559.92 ;
        LAYER Metal4 ;
        RECT  0.33 0.33 114.68 559.92 ;
        LAYER Metal5 ;
        RECT  114.65 0.33 114.68 559.92 ;
        RECT  103.70 2.20 114.65 559.92 ;
        RECT  4.05 2.20 14.70 559.92 ;
        RECT  2.20 0.33 4.05 559.92 ;
        RECT  0.33 0.33 2.20 59.75 ;
        RECT  0.33 108.90 2.20 109.60 ;
        RECT  0.33 241.90 2.20 242.60 ;
        RECT  0.33 380.90 2.20 559.92 ;
        RECT  14.70 0.33 103.70 559.92 ;
    END
END iobuf3_16pu_8

MACRO iobufdv_16_12
    CLASS PAD ;
    FOREIGN iobufdv_16_12  0.00 -38.75 N  ;
    ORIGIN 0.00 39.15 ;
    SIZE 115.00 BY 600.00 ;
    SYMMETRY x y r90 ;
    SITE io_site ;
     PIN en USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  60.95 -0.40 61.55 0.30 ;
        END
    END en
    PIN pad USE SIGNAL ; DIRECTION INOUT ;
        PORT
        LAYER Metal3 ;
        RECT  3.00 383.00 112.00 544.25 ;
        END
    END pad
    PIN do USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  25.95 -0.40 26.55 0.30 ;
        END
    END do
    PIN di  USE SIGNAL ; DIRECTION OUTPUT ;
        PORT
        LAYER Metal1 ;
        RECT  87.15 -0.40 87.75 0.30 ;
        END
    END di
    PIN vdd!
        USE power ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        LAYER Metal3 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        END
    END vdd!
    PIN vss!
        USE ground ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        LAYER Metal3 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        END
    END vss!
    OBS
        LAYER Metal1 ;
        RECT  88.35 -0.40 114.75 560.00 ;
        RECT  86.55 0.90 88.35 560.00 ;
        RECT  62.15 -0.40 86.55 560.00 ;
        RECT  60.35 0.90 62.15 560.00 ;
        RECT  27.15 -0.40 60.35 560.00 ;
        RECT  25.35 0.90 27.15 560.00 ;
        RECT  0.25 -0.40 25.35 560.00 ;
        LAYER Metal2 ;
        RECT  0.33 0.33 114.68 559.92 ;
        LAYER Metal3 ;
        RECT  114.65 0.33 114.68 559.92 ;
        RECT  103.70 2.20 114.65 559.92 ;
        RECT  4.05 2.20 14.70 559.92 ;
        RECT  2.20 0.33 4.05 559.92 ;
        RECT  0.33 0.33 2.20 59.75 ;
        RECT  0.33 108.90 2.20 109.60 ;
        RECT  0.33 241.90 2.20 242.60 ;
        RECT  0.33 380.90 2.20 559.92 ;
        RECT  14.70 0.33 103.70 559.92 ;
    END
END iobufdv_16_12

MACRO iobufdv_16_4
    CLASS PAD ;
    FOREIGN iobufdv_16_4  0.00 -38.75 N  ;
    ORIGIN 0.00 39.15 ;
    SIZE 115.00 BY 600.00 ;
    SYMMETRY x y r90 ;
    SITE io_site ;
     PIN en USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  60.95 -0.40 61.55 0.30 ;
        END
    END en
    PIN pad USE SIGNAL ; DIRECTION INOUT ;
        PORT
        LAYER Metal3 ;
        RECT  3.00 383.00 112.00 544.25 ;
        END
    END pad
    PIN do USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  25.95 -0.40 26.55 0.30 ;
        END
    END do
    PIN di  USE SIGNAL ; DIRECTION OUTPUT ;
        PORT
        LAYER Metal1 ;
        RECT  87.15 -0.40 87.75 0.30 ;
        END
    END di
    PIN vdd!
        USE power ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        LAYER Metal3 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        END
    END vdd!
    PIN vss!
        USE ground ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        LAYER Metal3 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        END
    END vss!
    OBS
        LAYER Metal1 ;
        RECT  88.35 -0.40 114.75 560.00 ;
        RECT  86.55 0.90 88.35 560.00 ;
        RECT  62.15 -0.40 86.55 560.00 ;
        RECT  60.35 0.90 62.15 560.00 ;
        RECT  27.15 -0.40 60.35 560.00 ;
        RECT  25.35 0.90 27.15 560.00 ;
        RECT  0.25 -0.40 25.35 560.00 ;
        LAYER Metal2 ;
        RECT  0.33 0.33 114.68 559.92 ;
        LAYER Metal3 ;
        RECT  114.65 0.33 114.68 559.92 ;
        RECT  103.70 2.20 114.65 559.92 ;
        RECT  4.05 2.20 14.70 559.92 ;
        RECT  2.20 0.33 4.05 559.92 ;
        RECT  0.33 0.33 2.20 59.75 ;
        RECT  0.33 108.90 2.20 109.60 ;
        RECT  0.33 241.90 2.20 242.60 ;
        RECT  0.33 380.90 2.20 559.92 ;
        RECT  14.70 0.33 103.70 559.92 ;
    END
END iobufdv_16_4

MACRO iobufdv_16_8
    CLASS PAD ;
    FOREIGN iobufdv_16_8  0.00 -38.75 N  ;
    ORIGIN 0.00 39.15 ;
    SIZE 115.00 BY 600.00 ;
    SYMMETRY x y r90 ;
    SITE io_site ;
     PIN en USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  60.95 -0.40 61.55 0.30 ;
        END
    END en
    PIN pad USE SIGNAL ; DIRECTION INOUT ;
        PORT
        LAYER Metal3 ;
        RECT  3.00 383.00 112.00 544.25 ;
        END
    END pad
    PIN do USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  25.95 -0.40 26.55 0.30 ;
        END
    END do
    PIN di  USE SIGNAL ; DIRECTION OUTPUT ;
        PORT
        LAYER Metal1 ;
        RECT  87.15 -0.40 87.75 0.30 ;
        END
    END di
    PIN vdd!
        USE power ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        LAYER Metal3 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        END
    END vdd!
    PIN vss!
        USE ground ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        LAYER Metal3 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        END
    END vss!
    OBS
        LAYER Metal1 ;
        RECT  88.35 -0.40 114.75 560.00 ;
        RECT  86.55 0.90 88.35 560.00 ;
        RECT  62.15 -0.40 86.55 560.00 ;
        RECT  60.35 0.90 62.15 560.00 ;
        RECT  27.15 -0.40 60.35 560.00 ;
        RECT  25.35 0.90 27.15 560.00 ;
        RECT  0.25 -0.40 25.35 560.00 ;
        LAYER Metal2 ;
        RECT  0.33 0.33 114.68 559.92 ;
        LAYER Metal3 ;
        RECT  114.65 0.33 114.68 559.92 ;
        RECT  103.70 2.20 114.65 559.92 ;
        RECT  4.05 2.20 14.70 559.92 ;
        RECT  2.20 0.33 4.05 559.92 ;
        RECT  0.33 0.33 2.20 59.75 ;
        RECT  0.33 108.90 2.20 109.60 ;
        RECT  0.33 241.90 2.20 242.60 ;
        RECT  0.33 380.90 2.20 559.92 ;
        RECT  14.70 0.33 103.70 559.92 ;
    END
END iobufdv_16_8

MACRO iobufdv_16pd_12
    CLASS PAD ;
    FOREIGN iobufdv_16pd_12  0.00 -38.75 N  ;
    ORIGIN 0.00 39.15 ;
    SIZE 115.00 BY 600.00 ;
    SYMMETRY x y r90 ;
    SITE io_site ;
     PIN en USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  60.95 -0.40 61.55 0.30 ;
        END
    END en
    PIN pad USE SIGNAL ; DIRECTION INOUT ;
        PORT
        LAYER Metal3 ;
        RECT  3.00 383.00 112.00 544.25 ;
        END
    END pad
    PIN do USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  25.95 -0.40 26.55 0.30 ;
        END
    END do
    PIN di  USE SIGNAL ; DIRECTION OUTPUT ;
        PORT
        LAYER Metal1 ;
        RECT  87.15 -0.40 87.75 0.30 ;
        END
    END di
    PIN vdd!
        USE power ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        LAYER Metal3 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        END
    END vdd!
    PIN vss!
        USE ground ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        LAYER Metal3 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        END
    END vss!
    OBS
        LAYER Metal1 ;
        RECT  88.35 -0.40 114.75 560.00 ;
        RECT  86.55 0.90 88.35 560.00 ;
        RECT  62.15 -0.40 86.55 560.00 ;
        RECT  60.35 0.90 62.15 560.00 ;
        RECT  27.15 -0.40 60.35 560.00 ;
        RECT  25.35 0.90 27.15 560.00 ;
        RECT  0.25 -0.40 25.35 560.00 ;
        LAYER Metal2 ;
        RECT  0.33 0.33 114.68 559.92 ;
        LAYER Metal3 ;
        RECT  114.65 0.33 114.68 559.92 ;
        RECT  103.70 2.20 114.65 559.92 ;
        RECT  4.05 2.20 14.70 559.92 ;
        RECT  2.20 0.33 4.05 559.92 ;
        RECT  0.33 0.33 2.20 59.75 ;
        RECT  0.33 108.90 2.20 109.60 ;
        RECT  0.33 241.90 2.20 242.60 ;
        RECT  0.33 380.90 2.20 559.92 ;
        RECT  14.70 0.33 103.70 559.92 ;
    END
END iobufdv_16pd_12

MACRO iobufdv_16pd_4
    CLASS PAD ;
    FOREIGN iobufdv_16pd_4  0.00 -38.75 N  ;
    ORIGIN 0.00 39.15 ;
    SIZE 115.00 BY 600.00 ;
    SYMMETRY x y r90 ;
    SITE io_site ;
     PIN en USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  60.95 -0.40 61.55 0.30 ;
        END
    END en
    PIN pad USE SIGNAL ; DIRECTION INOUT ;
        PORT
        LAYER Metal3 ;
        RECT  3.00 383.00 112.00 544.25 ;
        END
    END pad
    PIN do USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  25.95 -0.40 26.55 0.30 ;
        END
    END do
    PIN di  USE SIGNAL ; DIRECTION OUTPUT ;
        PORT
        LAYER Metal1 ;
        RECT  87.15 -0.40 87.75 0.30 ;
        END
    END di
    PIN vdd!
        USE power ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        LAYER Metal3 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        END
    END vdd!
    PIN vss!
        USE ground ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        LAYER Metal3 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        END
    END vss!
    OBS
        LAYER Metal1 ;
        RECT  88.35 -0.40 114.75 560.00 ;
        RECT  86.55 0.90 88.35 560.00 ;
        RECT  62.15 -0.40 86.55 560.00 ;
        RECT  60.35 0.90 62.15 560.00 ;
        RECT  27.15 -0.40 60.35 560.00 ;
        RECT  25.35 0.90 27.15 560.00 ;
        RECT  0.25 -0.40 25.35 560.00 ;
        LAYER Metal2 ;
        RECT  0.33 0.33 114.68 559.92 ;
        LAYER Metal3 ;
        RECT  114.65 0.33 114.68 559.92 ;
        RECT  103.70 2.20 114.65 559.92 ;
        RECT  4.05 2.20 14.70 559.92 ;
        RECT  2.20 0.33 4.05 559.92 ;
        RECT  0.33 0.33 2.20 59.75 ;
        RECT  0.33 108.90 2.20 109.60 ;
        RECT  0.33 241.90 2.20 242.60 ;
        RECT  0.33 380.90 2.20 559.92 ;
        RECT  14.70 0.33 103.70 559.92 ;
    END
END iobufdv_16pd_4

MACRO iobufdv_16pd_8
    CLASS PAD ;
    FOREIGN iobufdv_16pd_8  0.00 -38.75 N  ;
    ORIGIN 0.00 39.15 ;
    SIZE 115.00 BY 600.00 ;
    SYMMETRY x y r90 ;
    SITE io_site ;
     PIN en USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  60.95 -0.40 61.55 0.30 ;
        END
    END en
    PIN pad USE SIGNAL ; DIRECTION INOUT ;
        PORT
        LAYER Metal3 ;
        RECT  3.00 383.00 112.00 544.25 ;
        END
    END pad
    PIN do USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  25.95 -0.40 26.55 0.30 ;
        END
    END do
    PIN di  USE SIGNAL ; DIRECTION OUTPUT ;
        PORT
        LAYER Metal1 ;
        RECT  87.15 -0.40 87.75 0.30 ;
        END
    END di
    PIN vdd!
        USE power ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        LAYER Metal3 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        END
    END vdd!
    PIN vss!
        USE ground ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        LAYER Metal3 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        END
    END vss!
    OBS
        LAYER Metal1 ;
        RECT  88.35 -0.40 114.75 560.00 ;
        RECT  86.55 0.90 88.35 560.00 ;
        RECT  62.15 -0.40 86.55 560.00 ;
        RECT  60.35 0.90 62.15 560.00 ;
        RECT  27.15 -0.40 60.35 560.00 ;
        RECT  25.35 0.90 27.15 560.00 ;
        RECT  0.25 -0.40 25.35 560.00 ;
        LAYER Metal2 ;
        RECT  0.33 0.33 114.68 559.92 ;
        LAYER Metal3 ;
        RECT  114.65 0.33 114.68 559.92 ;
        RECT  103.70 2.20 114.65 559.92 ;
        RECT  4.05 2.20 14.70 559.92 ;
        RECT  2.20 0.33 4.05 559.92 ;
        RECT  0.33 0.33 2.20 59.75 ;
        RECT  0.33 108.90 2.20 109.60 ;
        RECT  0.33 241.90 2.20 242.60 ;
        RECT  0.33 380.90 2.20 559.92 ;
        RECT  14.70 0.33 103.70 559.92 ;
    END
END iobufdv_16pd_8

MACRO iobufdv_16pu_12
    CLASS PAD ;
    FOREIGN iobufdv_16pu_12  0.00 -38.75 N  ;
    ORIGIN 0.00 39.15 ;
    SIZE 115.00 BY 600.00 ;
    SYMMETRY x y r90 ;
    SITE io_site ;
     PIN en USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  60.95 -0.40 61.55 0.30 ;
        END
    END en
    PIN pad USE SIGNAL ; DIRECTION INOUT ;
        PORT
        LAYER Metal3 ;
        RECT  3.00 383.00 112.00 544.25 ;
        END
    END pad
    PIN do USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  25.95 -0.40 26.55 0.30 ;
        END
    END do
    PIN di  USE SIGNAL ; DIRECTION OUTPUT ;
        PORT
        LAYER Metal1 ;
        RECT  87.15 -0.40 87.75 0.30 ;
        END
    END di
    PIN vdd!
        USE power ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        LAYER Metal3 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        END
    END vdd!
    PIN vss!
        USE ground ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        LAYER Metal3 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        END
    END vss!
    OBS
        LAYER Metal1 ;
        RECT  88.35 -0.40 114.75 560.00 ;
        RECT  86.55 0.90 88.35 560.00 ;
        RECT  62.15 -0.40 86.55 560.00 ;
        RECT  60.35 0.90 62.15 560.00 ;
        RECT  27.15 -0.40 60.35 560.00 ;
        RECT  25.35 0.90 27.15 560.00 ;
        RECT  0.25 -0.40 25.35 560.00 ;
        LAYER Metal2 ;
        RECT  0.33 0.33 114.68 559.92 ;
        LAYER Metal3 ;
        RECT  114.65 0.33 114.68 559.92 ;
        RECT  103.70 2.20 114.65 559.92 ;
        RECT  4.05 2.20 14.70 559.92 ;
        RECT  2.20 0.33 4.05 559.92 ;
        RECT  0.33 0.33 2.20 59.75 ;
        RECT  0.33 108.90 2.20 109.60 ;
        RECT  0.33 241.90 2.20 242.60 ;
        RECT  0.33 380.90 2.20 559.92 ;
        RECT  14.70 0.33 103.70 559.92 ;
    END
END iobufdv_16pu_12

MACRO iobufdv_16pu_4
    CLASS PAD ;
    FOREIGN iobufdv_16pu_4  0.00 -38.75 N  ;
    ORIGIN 0.00 39.15 ;
    SIZE 115.00 BY 600.00 ;
    SYMMETRY x y r90 ;
    SITE io_site ;
     PIN en USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  60.95 -0.40 61.55 0.30 ;
        END
    END en
    PIN pad USE SIGNAL ; DIRECTION INOUT ;
        PORT
        LAYER Metal3 ;
        RECT  3.00 383.00 112.00 544.25 ;
        END
    END pad
    PIN do USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  25.95 -0.40 26.55 0.30 ;
        END
    END do
    PIN di  USE SIGNAL ; DIRECTION OUTPUT ;
        PORT
        LAYER Metal1 ;
        RECT  87.15 -0.40 87.75 0.30 ;
        END
    END di
    PIN vdd!
        USE power ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        LAYER Metal3 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        END
    END vdd!
    PIN vss!
        USE ground ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        LAYER Metal3 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        END
    END vss!
    OBS
        LAYER Metal1 ;
        RECT  88.35 -0.40 114.75 560.00 ;
        RECT  86.55 0.90 88.35 560.00 ;
        RECT  62.15 -0.40 86.55 560.00 ;
        RECT  60.35 0.90 62.15 560.00 ;
        RECT  27.15 -0.40 60.35 560.00 ;
        RECT  25.35 0.90 27.15 560.00 ;
        RECT  0.25 -0.40 25.35 560.00 ;
        LAYER Metal2 ;
        RECT  0.33 0.33 114.68 559.92 ;
        LAYER Metal3 ;
        RECT  114.65 0.33 114.68 559.92 ;
        RECT  103.70 2.20 114.65 559.92 ;
        RECT  4.05 2.20 14.70 559.92 ;
        RECT  2.20 0.33 4.05 559.92 ;
        RECT  0.33 0.33 2.20 59.75 ;
        RECT  0.33 108.90 2.20 109.60 ;
        RECT  0.33 241.90 2.20 242.60 ;
        RECT  0.33 380.90 2.20 559.92 ;
        RECT  14.70 0.33 103.70 559.92 ;
    END
END iobufdv_16pu_4

MACRO iobufdv_16pu_8
    CLASS PAD ;
    FOREIGN iobufdv_16pu_8  0.00 -38.75 N  ;
    ORIGIN 0.00 39.15 ;
    SIZE 115.00 BY 600.00 ;
    SYMMETRY x y r90 ;
    SITE io_site ;
     PIN en USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  60.95 -0.40 61.55 0.30 ;
        END
    END en
    PIN pad USE SIGNAL ; DIRECTION INOUT ;
        PORT
        LAYER Metal3 ;
        RECT  3.00 383.00 112.00 544.25 ;
        END
    END pad
    PIN do USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  25.95 -0.40 26.55 0.30 ;
        END
    END do
    PIN di  USE SIGNAL ; DIRECTION OUTPUT ;
        PORT
        LAYER Metal1 ;
        RECT  87.15 -0.40 87.75 0.30 ;
        END
    END di
    PIN vdd!
        USE power ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        LAYER Metal3 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        END
    END vdd!
    PIN vss!
        USE ground ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        LAYER Metal3 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        END
    END vss!
    OBS
        LAYER Metal1 ;
        RECT  88.35 -0.40 114.75 560.00 ;
        RECT  86.55 0.90 88.35 560.00 ;
        RECT  62.15 -0.40 86.55 560.00 ;
        RECT  60.35 0.90 62.15 560.00 ;
        RECT  27.15 -0.40 60.35 560.00 ;
        RECT  25.35 0.90 27.15 560.00 ;
        RECT  0.25 -0.40 25.35 560.00 ;
        LAYER Metal2 ;
        RECT  0.33 0.33 114.68 559.92 ;
        LAYER Metal3 ;
        RECT  114.65 0.33 114.68 559.92 ;
        RECT  103.70 2.20 114.65 559.92 ;
        RECT  4.05 2.20 14.70 559.92 ;
        RECT  2.20 0.33 4.05 559.92 ;
        RECT  0.33 0.33 2.20 59.75 ;
        RECT  0.33 108.90 2.20 109.60 ;
        RECT  0.33 241.90 2.20 242.60 ;
        RECT  0.33 380.90 2.20 559.92 ;
        RECT  14.70 0.33 103.70 559.92 ;
    END
END iobufdv_16pu_8

MACRO iobufs2_16_12
    CLASS PAD ;
    FOREIGN iobufs2_16_12  0.00 -38.75 N  ;
    ORIGIN 0.00 39.15 ;
    SIZE 115.00 BY 600.00 ;
    SYMMETRY x y r90 ;
    SITE io_site ;
     PIN en USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  60.95 -0.40 61.55 0.30 ;
        END
    END en
    PIN pad USE SIGNAL ; DIRECTION INOUT ;
        PORT
        LAYER Metal3 ;
        RECT  3.00 383.00 112.00 544.25 ;
        END
    END pad
    PIN do USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  25.95 -0.40 26.55 0.30 ;
        END
    END do
    PIN di  USE SIGNAL ; DIRECTION OUTPUT ;
        PORT
        LAYER Metal1 ;
        RECT  87.15 -0.40 87.75 0.30 ;
        END
    END di
    PIN vdd!
        USE power ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        LAYER Metal3 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        END
    END vdd!
    PIN vss!
        USE ground ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        LAYER Metal3 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        END
    END vss!
    OBS
        LAYER Metal1 ;
        RECT  88.35 -0.40 114.75 560.00 ;
        RECT  86.55 0.90 88.35 560.00 ;
        RECT  62.15 -0.40 86.55 560.00 ;
        RECT  60.35 0.90 62.15 560.00 ;
        RECT  27.15 -0.40 60.35 560.00 ;
        RECT  25.35 0.90 27.15 560.00 ;
        RECT  0.25 -0.40 25.35 560.00 ;
        LAYER Metal2 ;
        RECT  0.33 0.33 114.68 559.92 ;
        LAYER Metal3 ;
        RECT  114.65 0.33 114.68 559.92 ;
        RECT  103.70 2.20 114.65 559.92 ;
        RECT  4.05 2.20 14.70 559.92 ;
        RECT  2.20 0.33 4.05 559.92 ;
        RECT  0.33 0.33 2.20 59.75 ;
        RECT  0.33 108.90 2.20 109.60 ;
        RECT  0.33 241.90 2.20 242.60 ;
        RECT  0.33 380.90 2.20 559.92 ;
        RECT  14.70 0.33 103.70 559.92 ;
    END
END iobufs2_16_12

MACRO iobufs2_16_4
    CLASS PAD ;
    FOREIGN iobufs2_16_4  0.00 -38.75 N  ;
    ORIGIN 0.00 39.15 ;
    SIZE 115.00 BY 600.00 ;
    SYMMETRY x y r90 ;
    SITE io_site ;
     PIN en USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  60.95 -0.40 61.55 0.30 ;
        END
    END en
    PIN pad USE SIGNAL ; DIRECTION INOUT ;
        PORT
        LAYER Metal3 ;
        RECT  3.00 383.00 112.00 544.25 ;
        END
    END pad
    PIN do USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  25.95 -0.40 26.55 0.30 ;
        END
    END do
    PIN di  USE SIGNAL ; DIRECTION OUTPUT ;
        PORT
        LAYER Metal1 ;
        RECT  87.15 -0.40 87.75 0.30 ;
        END
    END di
    PIN vdd!
        USE power ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        LAYER Metal3 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        END
    END vdd!
    PIN vss!
        USE ground ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        LAYER Metal3 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        END
    END vss!
    OBS
        LAYER Metal1 ;
        RECT  88.35 -0.40 114.75 560.00 ;
        RECT  86.55 0.90 88.35 560.00 ;
        RECT  62.15 -0.40 86.55 560.00 ;
        RECT  60.35 0.90 62.15 560.00 ;
        RECT  27.15 -0.40 60.35 560.00 ;
        RECT  25.35 0.90 27.15 560.00 ;
        RECT  0.25 -0.40 25.35 560.00 ;
        LAYER Metal2 ;
        RECT  0.33 0.33 114.68 559.92 ;
        LAYER Metal3 ;
        RECT  114.65 0.33 114.68 559.92 ;
        RECT  103.70 2.20 114.65 559.92 ;
        RECT  4.05 2.20 14.70 559.92 ;
        RECT  2.20 0.33 4.05 559.92 ;
        RECT  0.33 0.33 2.20 59.75 ;
        RECT  0.33 108.90 2.20 109.60 ;
        RECT  0.33 241.90 2.20 242.60 ;
        RECT  0.33 380.90 2.20 559.92 ;
        RECT  14.70 0.33 103.70 559.92 ;
    END
END iobufs2_16_4

MACRO iobufs2_16_8
    CLASS PAD ;
    FOREIGN iobufs2_16_8  0.00 -38.75 N  ;
    ORIGIN 0.00 39.15 ;
    SIZE 115.00 BY 600.00 ;
    SYMMETRY x y r90 ;
    SITE io_site ;
     PIN en USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  60.95 -0.40 61.55 0.30 ;
        END
    END en
    PIN pad USE SIGNAL ; DIRECTION INOUT ;
        PORT
        LAYER Metal3 ;
        RECT  3.00 383.00 112.00 544.25 ;
        END
    END pad
    PIN do USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  25.95 -0.40 26.55 0.30 ;
        END
    END do
    PIN di  USE SIGNAL ; DIRECTION OUTPUT ;
        PORT
        LAYER Metal1 ;
        RECT  87.15 -0.40 87.75 0.30 ;
        END
    END di
    PIN vdd!
        USE power ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        LAYER Metal3 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        END
    END vdd!
    PIN vss!
        USE ground ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        LAYER Metal3 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        END
    END vss!
    OBS
        LAYER Metal1 ;
        RECT  88.35 -0.40 114.75 560.00 ;
        RECT  86.55 0.90 88.35 560.00 ;
        RECT  62.15 -0.40 86.55 560.00 ;
        RECT  60.35 0.90 62.15 560.00 ;
        RECT  27.15 -0.40 60.35 560.00 ;
        RECT  25.35 0.90 27.15 560.00 ;
        RECT  0.25 -0.40 25.35 560.00 ;
        LAYER Metal2 ;
        RECT  0.33 0.33 114.68 559.92 ;
        LAYER Metal3 ;
        RECT  114.65 0.33 114.68 559.92 ;
        RECT  103.70 2.20 114.65 559.92 ;
        RECT  4.05 2.20 14.70 559.92 ;
        RECT  2.20 0.33 4.05 559.92 ;
        RECT  0.33 0.33 2.20 59.75 ;
        RECT  0.33 108.90 2.20 109.60 ;
        RECT  0.33 241.90 2.20 242.60 ;
        RECT  0.33 380.90 2.20 559.92 ;
        RECT  14.70 0.33 103.70 559.92 ;
    END
END iobufs2_16_8

MACRO iobufs2_16pd_12
    CLASS PAD ;
    FOREIGN iobufs2_16pd_12  0.00 -38.75 N  ;
    ORIGIN 0.00 39.15 ;
    SIZE 115.00 BY 600.00 ;
    SYMMETRY x y r90 ;
    SITE io_site ;
     PIN en USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  60.95 -0.40 61.55 0.30 ;
        END
    END en
    PIN pad USE SIGNAL ; DIRECTION INOUT ;
        PORT
        LAYER Metal3 ;
        RECT  3.00 383.00 112.00 544.25 ;
        END
    END pad
    PIN do USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  25.95 -0.40 26.55 0.30 ;
        END
    END do
    PIN di  USE SIGNAL ; DIRECTION OUTPUT ;
        PORT
        LAYER Metal1 ;
        RECT  87.15 -0.40 87.75 0.30 ;
        END
    END di
    PIN vdd!
        USE power ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        LAYER Metal3 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        END
    END vdd!
    PIN vss!
        USE ground ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        LAYER Metal3 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        END
    END vss!
    OBS
        LAYER Metal1 ;
        RECT  88.35 -0.40 114.75 560.00 ;
        RECT  86.55 0.90 88.35 560.00 ;
        RECT  62.15 -0.40 86.55 560.00 ;
        RECT  60.35 0.90 62.15 560.00 ;
        RECT  27.15 -0.40 60.35 560.00 ;
        RECT  25.35 0.90 27.15 560.00 ;
        RECT  0.25 -0.40 25.35 560.00 ;
        LAYER Metal2 ;
        RECT  0.33 0.33 114.68 559.92 ;
        LAYER Metal3 ;
        RECT  114.65 0.33 114.68 559.92 ;
        RECT  103.70 2.20 114.65 559.92 ;
        RECT  4.05 2.20 14.70 559.92 ;
        RECT  2.20 0.33 4.05 559.92 ;
        RECT  0.33 0.33 2.20 59.75 ;
        RECT  0.33 108.90 2.20 109.60 ;
        RECT  0.33 241.90 2.20 242.60 ;
        RECT  0.33 380.90 2.20 559.92 ;
        RECT  14.70 0.33 103.70 559.92 ;
    END
END iobufs2_16pd_12

MACRO iobufs2_16pd_4
    CLASS PAD ;
    FOREIGN iobufs2_16pd_4  0.00 -38.75 N  ;
    ORIGIN 0.00 39.15 ;
    SIZE 115.00 BY 600.00 ;
    SYMMETRY x y r90 ;
    SITE io_site ;
     PIN en USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  60.95 -0.40 61.55 0.30 ;
        END
    END en
    PIN pad USE SIGNAL ; DIRECTION INOUT ;
        PORT
        LAYER Metal3 ;
        RECT  3.00 383.00 112.00 544.25 ;
        END
    END pad
    PIN do USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  25.95 -0.40 26.55 0.30 ;
        END
    END do
    PIN di  USE SIGNAL ; DIRECTION OUTPUT ;
        PORT
        LAYER Metal1 ;
        RECT  87.15 -0.40 87.75 0.30 ;
        END
    END di
    PIN vdd!
        USE power ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        LAYER Metal3 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        END
    END vdd!
    PIN vss!
        USE ground ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        LAYER Metal3 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        END
    END vss!
    OBS
        LAYER Metal1 ;
        RECT  88.35 -0.40 114.75 560.00 ;
        RECT  86.55 0.90 88.35 560.00 ;
        RECT  62.15 -0.40 86.55 560.00 ;
        RECT  60.35 0.90 62.15 560.00 ;
        RECT  27.15 -0.40 60.35 560.00 ;
        RECT  25.35 0.90 27.15 560.00 ;
        RECT  0.25 -0.40 25.35 560.00 ;
        LAYER Metal2 ;
        RECT  0.33 0.33 114.68 559.92 ;
        LAYER Metal3 ;
        RECT  114.65 0.33 114.68 559.92 ;
        RECT  103.70 2.20 114.65 559.92 ;
        RECT  4.05 2.20 14.70 559.92 ;
        RECT  2.20 0.33 4.05 559.92 ;
        RECT  0.33 0.33 2.20 59.75 ;
        RECT  0.33 108.90 2.20 109.60 ;
        RECT  0.33 241.90 2.20 242.60 ;
        RECT  0.33 380.90 2.20 559.92 ;
        RECT  14.70 0.33 103.70 559.92 ;
    END
END iobufs2_16pd_4

MACRO iobufs2_16pd_8
    CLASS PAD ;
    FOREIGN iobufs2_16pd_8  0.00 -38.75 N  ;
    ORIGIN 0.00 39.15 ;
    SIZE 115.00 BY 600.00 ;
    SYMMETRY x y r90 ;
    SITE io_site ;
     PIN en USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  60.95 -0.40 61.55 0.30 ;
        END
    END en
    PIN pad USE SIGNAL ; DIRECTION INOUT ;
        PORT
        LAYER Metal3 ;
        RECT  3.00 383.00 112.00 544.25 ;
        END
    END pad
    PIN do USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  25.95 -0.40 26.55 0.30 ;
        END
    END do
    PIN di  USE SIGNAL ; DIRECTION OUTPUT ;
        PORT
        LAYER Metal1 ;
        RECT  87.15 -0.40 87.75 0.30 ;
        END
    END di
    PIN vdd!
        USE power ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        LAYER Metal3 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        END
    END vdd!
    PIN vss!
        USE ground ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        LAYER Metal3 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        END
    END vss!
    OBS
        LAYER Metal1 ;
        RECT  88.35 -0.40 114.75 560.00 ;
        RECT  86.55 0.90 88.35 560.00 ;
        RECT  62.15 -0.40 86.55 560.00 ;
        RECT  60.35 0.90 62.15 560.00 ;
        RECT  27.15 -0.40 60.35 560.00 ;
        RECT  25.35 0.90 27.15 560.00 ;
        RECT  0.25 -0.40 25.35 560.00 ;
        LAYER Metal2 ;
        RECT  0.33 0.33 114.68 559.92 ;
        LAYER Metal3 ;
        RECT  114.65 0.33 114.68 559.92 ;
        RECT  103.70 2.20 114.65 559.92 ;
        RECT  4.05 2.20 14.70 559.92 ;
        RECT  2.20 0.33 4.05 559.92 ;
        RECT  0.33 0.33 2.20 59.75 ;
        RECT  0.33 108.90 2.20 109.60 ;
        RECT  0.33 241.90 2.20 242.60 ;
        RECT  0.33 380.90 2.20 559.92 ;
        RECT  14.70 0.33 103.70 559.92 ;
    END
END iobufs2_16pd_8

MACRO iobufs2_16pu_12
    CLASS PAD ;
    FOREIGN iobufs2_16pu_12  0.00 -38.75 N  ;
    ORIGIN 0.00 39.15 ;
    SIZE 115.00 BY 600.00 ;
    SYMMETRY x y r90 ;
    SITE io_site ;
     PIN en USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  60.95 -0.40 61.55 0.30 ;
        END
    END en
    PIN pad USE SIGNAL ; DIRECTION INOUT ;
        PORT
        LAYER Metal3 ;
        RECT  3.00 383.00 112.00 544.25 ;
        END
    END pad
    PIN do USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  25.95 -0.40 26.55 0.30 ;
        END
    END do
    PIN di  USE SIGNAL ; DIRECTION OUTPUT ;
        PORT
        LAYER Metal1 ;
        RECT  87.15 -0.40 87.75 0.30 ;
        END
    END di
    PIN vdd!
        USE power ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        LAYER Metal3 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        END
    END vdd!
    PIN vss!
        USE ground ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        LAYER Metal3 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        END
    END vss!
    OBS
        LAYER Metal1 ;
        RECT  88.35 -0.40 114.75 560.00 ;
        RECT  86.55 0.90 88.35 560.00 ;
        RECT  62.15 -0.40 86.55 560.00 ;
        RECT  60.35 0.90 62.15 560.00 ;
        RECT  27.15 -0.40 60.35 560.00 ;
        RECT  25.35 0.90 27.15 560.00 ;
        RECT  0.25 -0.40 25.35 560.00 ;
        LAYER Metal2 ;
        RECT  0.33 0.33 114.68 559.92 ;
        LAYER Metal3 ;
        RECT  114.65 0.33 114.68 559.92 ;
        RECT  103.70 2.20 114.65 559.92 ;
        RECT  4.05 2.20 14.70 559.92 ;
        RECT  2.20 0.33 4.05 559.92 ;
        RECT  0.33 0.33 2.20 59.75 ;
        RECT  0.33 108.90 2.20 109.60 ;
        RECT  0.33 241.90 2.20 242.60 ;
        RECT  0.33 380.90 2.20 559.92 ;
        RECT  14.70 0.33 103.70 559.92 ;
    END
END iobufs2_16pu_12

MACRO iobufs2_16pu_4
    CLASS PAD ;
    FOREIGN iobufs2_16pu_4  0.00 -38.75 N  ;
    ORIGIN 0.00 39.15 ;
    SIZE 115.00 BY 600.00 ;
    SYMMETRY x y r90 ;
    SITE io_site ;
     PIN en USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  60.95 -0.40 61.55 0.30 ;
        END
    END en
    PIN pad USE SIGNAL ; DIRECTION INOUT ;
        PORT
        LAYER Metal3 ;
        RECT  3.00 383.00 112.00 544.25 ;
        END
    END pad
    PIN do USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  25.95 -0.40 26.55 0.30 ;
        END
    END do
    PIN di  USE SIGNAL ; DIRECTION OUTPUT ;
        PORT
        LAYER Metal1 ;
        RECT  87.15 -0.40 87.75 0.30 ;
        END
    END di
    PIN vdd!
        USE power ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        LAYER Metal3 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        END
    END vdd!
    PIN vss!
        USE ground ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        LAYER Metal3 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        END
    END vss!
    OBS
        LAYER Metal1 ;
        RECT  88.35 -0.40 114.75 560.00 ;
        RECT  86.55 0.90 88.35 560.00 ;
        RECT  62.15 -0.40 86.55 560.00 ;
        RECT  60.35 0.90 62.15 560.00 ;
        RECT  27.15 -0.40 60.35 560.00 ;
        RECT  25.35 0.90 27.15 560.00 ;
        RECT  0.25 -0.40 25.35 560.00 ;
        LAYER Metal2 ;
        RECT  0.33 0.33 114.68 559.92 ;
        LAYER Metal3 ;
        RECT  114.65 0.33 114.68 559.92 ;
        RECT  103.70 2.20 114.65 559.92 ;
        RECT  4.05 2.20 14.70 559.92 ;
        RECT  2.20 0.33 4.05 559.92 ;
        RECT  0.33 0.33 2.20 59.75 ;
        RECT  0.33 108.90 2.20 109.60 ;
        RECT  0.33 241.90 2.20 242.60 ;
        RECT  0.33 380.90 2.20 559.92 ;
        RECT  14.70 0.33 103.70 559.92 ;
    END
END iobufs2_16pu_4

MACRO iobufs2_16pu_8
    CLASS PAD ;
    FOREIGN iobufs2_16pu_8  0.00 -38.75 N  ;
    ORIGIN 0.00 39.15 ;
    SIZE 115.00 BY 600.00 ;
    SYMMETRY x y r90 ;
    SITE io_site ;
     PIN en USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  60.95 -0.40 61.55 0.30 ;
        END
    END en
    PIN pad USE SIGNAL ; DIRECTION INOUT ;
        PORT
        LAYER Metal3 ;
        RECT  3.00 383.00 112.00 544.25 ;
        END
    END pad
    PIN do USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  25.95 -0.40 26.55 0.30 ;
        END
    END do
    PIN di  USE SIGNAL ; DIRECTION OUTPUT ;
        PORT
        LAYER Metal1 ;
        RECT  87.15 -0.40 87.75 0.30 ;
        END
    END di
    PIN vdd!
        USE power ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        LAYER Metal3 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        END
    END vdd!
    PIN vss!
        USE ground ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        LAYER Metal3 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        END
    END vss!
    OBS
        LAYER Metal1 ;
        RECT  88.35 -0.40 114.75 560.00 ;
        RECT  86.55 0.90 88.35 560.00 ;
        RECT  62.15 -0.40 86.55 560.00 ;
        RECT  60.35 0.90 62.15 560.00 ;
        RECT  27.15 -0.40 60.35 560.00 ;
        RECT  25.35 0.90 27.15 560.00 ;
        RECT  0.25 -0.40 25.35 560.00 ;
        LAYER Metal2 ;
        RECT  0.33 0.33 114.68 559.92 ;
        LAYER Metal3 ;
        RECT  114.65 0.33 114.68 559.92 ;
        RECT  103.70 2.20 114.65 559.92 ;
        RECT  4.05 2.20 14.70 559.92 ;
        RECT  2.20 0.33 4.05 559.92 ;
        RECT  0.33 0.33 2.20 59.75 ;
        RECT  0.33 108.90 2.20 109.60 ;
        RECT  0.33 241.90 2.20 242.60 ;
        RECT  0.33 380.90 2.20 559.92 ;
        RECT  14.70 0.33 103.70 559.92 ;
    END
END iobufs2_16pu_8

MACRO iobufs3_16_12
    CLASS PAD ;
    FOREIGN iobufs3_16_12  0.00 -38.75 N  ;
    ORIGIN 0.00 39.15 ;
    SIZE 115.00 BY 600.00 ;
    SYMMETRY x y r90 ;
    SITE io_site ;
     PIN en USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  60.95 -0.40 61.55 0.30 ;
        END
    END en
    PIN pad USE SIGNAL ; DIRECTION INOUT ;
        PORT
        LAYER Metal3 ;
        RECT  3.00 383.00 112.00 544.25 ;
        END
    END pad
    PIN do USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  25.95 -0.40 26.55 0.30 ;
        END
    END do
    PIN di  USE SIGNAL ; DIRECTION OUTPUT ;
        PORT
        LAYER Metal1 ;
        RECT  87.15 -0.40 87.75 0.30 ;
        END
    END di
    PIN vdd!
        USE power ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        LAYER Metal3 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        END
    END vdd!
    PIN vss!
        USE ground ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        LAYER Metal3 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        END
    END vss!
    OBS
        LAYER Metal1 ;
        RECT  88.35 -0.40 114.75 560.00 ;
        RECT  86.55 0.90 88.35 560.00 ;
        RECT  62.15 -0.40 86.55 560.00 ;
        RECT  60.35 0.90 62.15 560.00 ;
        RECT  27.15 -0.40 60.35 560.00 ;
        RECT  25.35 0.90 27.15 560.00 ;
        RECT  0.25 -0.40 25.35 560.00 ;
        LAYER Metal2 ;
        RECT  0.33 0.33 114.68 559.92 ;
        LAYER Metal3 ;
        RECT  114.65 0.33 114.68 559.92 ;
        RECT  103.70 2.20 114.65 559.92 ;
        RECT  4.05 2.20 14.70 559.92 ;
        RECT  2.20 0.33 4.05 559.92 ;
        RECT  0.33 0.33 2.20 59.75 ;
        RECT  0.33 108.90 2.20 109.60 ;
        RECT  0.33 241.90 2.20 242.60 ;
        RECT  0.33 380.90 2.20 559.92 ;
        RECT  14.70 0.33 103.70 559.92 ;
    END
END iobufs3_16_12

MACRO iobufs3_16_4
    CLASS PAD ;
    FOREIGN iobufs3_16_4  0.00 -38.75 N  ;
    ORIGIN 0.00 39.15 ;
    SIZE 115.00 BY 600.00 ;
    SYMMETRY x y r90 ;
    SITE io_site ;
     PIN en USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  60.95 -0.40 61.55 0.30 ;
        END
    END en
    PIN pad USE SIGNAL ; DIRECTION INOUT ;
        PORT
        LAYER Metal3 ;
        RECT  3.00 383.00 112.00 544.25 ;
        END
    END pad
    PIN do USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  25.95 -0.40 26.55 0.30 ;
        END
    END do
    PIN di  USE SIGNAL ; DIRECTION OUTPUT ;
        PORT
        LAYER Metal1 ;
        RECT  87.15 -0.40 87.75 0.30 ;
        END
    END di
    PIN vdd!
        USE power ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        LAYER Metal3 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        END
    END vdd!
    PIN vss!
        USE ground ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        LAYER Metal3 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        END
    END vss!
    OBS
        LAYER Metal1 ;
        RECT  88.35 -0.40 114.75 560.00 ;
        RECT  86.55 0.90 88.35 560.00 ;
        RECT  62.15 -0.40 86.55 560.00 ;
        RECT  60.35 0.90 62.15 560.00 ;
        RECT  27.15 -0.40 60.35 560.00 ;
        RECT  25.35 0.90 27.15 560.00 ;
        RECT  0.25 -0.40 25.35 560.00 ;
        LAYER Metal2 ;
        RECT  0.33 0.33 114.68 559.92 ;
        LAYER Metal3 ;
        RECT  114.65 0.33 114.68 559.92 ;
        RECT  103.70 2.20 114.65 559.92 ;
        RECT  4.05 2.20 14.70 559.92 ;
        RECT  2.20 0.33 4.05 559.92 ;
        RECT  0.33 0.33 2.20 59.75 ;
        RECT  0.33 108.90 2.20 109.60 ;
        RECT  0.33 241.90 2.20 242.60 ;
        RECT  0.33 380.90 2.20 559.92 ;
        RECT  14.70 0.33 103.70 559.92 ;
    END
END iobufs3_16_4

MACRO iobufs3_16_8
    CLASS PAD ;
    FOREIGN iobufs3_16_8  0.00 -38.75 N  ;
    ORIGIN 0.00 39.15 ;
    SIZE 115.00 BY 600.00 ;
    SYMMETRY x y r90 ;
    SITE io_site ;
     PIN en USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  60.95 -0.40 61.55 0.30 ;
        END
    END en
    PIN pad USE SIGNAL ; DIRECTION INOUT ;
        PORT
        LAYER Metal3 ;
        RECT  3.00 383.00 112.00 544.25 ;
        END
    END pad
    PIN do USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  25.95 -0.40 26.55 0.30 ;
        END
    END do
    PIN di  USE SIGNAL ; DIRECTION OUTPUT ;
        PORT
        LAYER Metal1 ;
        RECT  87.15 -0.40 87.75 0.30 ;
        END
    END di
    PIN vdd!
        USE power ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        LAYER Metal3 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        END
    END vdd!
    PIN vss!
        USE ground ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        LAYER Metal3 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        END
    END vss!
    OBS
        LAYER Metal1 ;
        RECT  88.35 -0.40 114.75 560.00 ;
        RECT  86.55 0.90 88.35 560.00 ;
        RECT  62.15 -0.40 86.55 560.00 ;
        RECT  60.35 0.90 62.15 560.00 ;
        RECT  27.15 -0.40 60.35 560.00 ;
        RECT  25.35 0.90 27.15 560.00 ;
        RECT  0.25 -0.40 25.35 560.00 ;
        LAYER Metal2 ;
        RECT  0.33 0.33 114.68 559.92 ;
        LAYER Metal3 ;
        RECT  114.65 0.33 114.68 559.92 ;
        RECT  103.70 2.20 114.65 559.92 ;
        RECT  4.05 2.20 14.70 559.92 ;
        RECT  2.20 0.33 4.05 559.92 ;
        RECT  0.33 0.33 2.20 59.75 ;
        RECT  0.33 108.90 2.20 109.60 ;
        RECT  0.33 241.90 2.20 242.60 ;
        RECT  0.33 380.90 2.20 559.92 ;
        RECT  14.70 0.33 103.70 559.92 ;
    END
END iobufs3_16_8

MACRO iobufs3_16pd_12
    CLASS PAD ;
    FOREIGN iobufs3_16pd_12  0.00 -38.75 N  ;
    ORIGIN 0.00 39.15 ;
    SIZE 115.00 BY 600.00 ;
    SYMMETRY x y r90 ;
    SITE io_site ;
     PIN en USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  60.95 -0.40 61.55 0.30 ;
        END
    END en
    PIN pad USE SIGNAL ; DIRECTION INOUT ;
        PORT
        LAYER Metal3 ;
        RECT  3.00 383.00 112.00 544.25 ;
        END
    END pad
    PIN do USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  25.95 -0.40 26.55 0.30 ;
        END
    END do
    PIN di  USE SIGNAL ; DIRECTION OUTPUT ;
        PORT
        LAYER Metal1 ;
        RECT  87.15 -0.40 87.75 0.30 ;
        END
    END di
    PIN vdd!
        USE power ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        LAYER Metal3 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        END
    END vdd!
    PIN vss!
        USE ground ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        LAYER Metal3 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        END
    END vss!
    OBS
        LAYER Metal1 ;
        RECT  88.35 -0.40 114.75 560.00 ;
        RECT  86.55 0.90 88.35 560.00 ;
        RECT  62.15 -0.40 86.55 560.00 ;
        RECT  60.35 0.90 62.15 560.00 ;
        RECT  27.15 -0.40 60.35 560.00 ;
        RECT  25.35 0.90 27.15 560.00 ;
        RECT  0.25 -0.40 25.35 560.00 ;
        LAYER Metal2 ;
        RECT  0.33 0.33 114.68 559.92 ;
        LAYER Metal3 ;
        RECT  114.65 0.33 114.68 559.92 ;
        RECT  103.70 2.20 114.65 559.92 ;
        RECT  4.05 2.20 14.70 559.92 ;
        RECT  2.20 0.33 4.05 559.92 ;
        RECT  0.33 0.33 2.20 59.75 ;
        RECT  0.33 108.90 2.20 109.60 ;
        RECT  0.33 241.90 2.20 242.60 ;
        RECT  0.33 380.90 2.20 559.92 ;
        RECT  14.70 0.33 103.70 559.92 ;
    END
END iobufs3_16pd_12

MACRO iobufs3_16pd_4
    CLASS PAD ;
    FOREIGN iobufs3_16pd_4  0.00 -38.75 N  ;
    ORIGIN 0.00 39.15 ;
    SIZE 115.00 BY 600.00 ;
    SYMMETRY x y r90 ;
    SITE io_site ;
     PIN en USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  60.95 -0.40 61.55 0.30 ;
        END
    END en
    PIN pad USE SIGNAL ; DIRECTION INOUT ;
        PORT
        LAYER Metal3 ;
        RECT  3.00 383.00 112.00 544.25 ;
        END
    END pad
    PIN do USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  25.95 -0.40 26.55 0.30 ;
        END
    END do
    PIN di  USE SIGNAL ; DIRECTION OUTPUT ;
        PORT
        LAYER Metal1 ;
        RECT  87.15 -0.40 87.75 0.30 ;
        END
    END di
    PIN vdd!
        USE power ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        LAYER Metal3 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        END
    END vdd!
    PIN vss!
        USE ground ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        LAYER Metal3 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        END
    END vss!
    OBS
        LAYER Metal1 ;
        RECT  88.35 -0.40 114.75 560.00 ;
        RECT  86.55 0.90 88.35 560.00 ;
        RECT  62.15 -0.40 86.55 560.00 ;
        RECT  60.35 0.90 62.15 560.00 ;
        RECT  27.15 -0.40 60.35 560.00 ;
        RECT  25.35 0.90 27.15 560.00 ;
        RECT  0.25 -0.40 25.35 560.00 ;
        LAYER Metal2 ;
        RECT  0.33 0.33 114.68 559.92 ;
        LAYER Metal3 ;
        RECT  114.65 0.33 114.68 559.92 ;
        RECT  103.70 2.20 114.65 559.92 ;
        RECT  4.05 2.20 14.70 559.92 ;
        RECT  2.20 0.33 4.05 559.92 ;
        RECT  0.33 0.33 2.20 59.75 ;
        RECT  0.33 108.90 2.20 109.60 ;
        RECT  0.33 241.90 2.20 242.60 ;
        RECT  0.33 380.90 2.20 559.92 ;
        RECT  14.70 0.33 103.70 559.92 ;
    END
END iobufs3_16pd_4

MACRO iobufs3_16pd_8
    CLASS PAD ;
    FOREIGN iobufs3_16pd_8  0.00 -38.75 N  ;
    ORIGIN 0.00 39.15 ;
    SIZE 115.00 BY 600.00 ;
    SYMMETRY x y r90 ;
    SITE io_site ;
     PIN en USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  60.95 -0.40 61.55 0.30 ;
        END
    END en
    PIN pad USE SIGNAL ; DIRECTION INOUT ;
        PORT
        LAYER Metal3 ;
        RECT  3.00 383.00 112.00 544.25 ;
        END
    END pad
    PIN do USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  25.95 -0.40 26.55 0.30 ;
        END
    END do
    PIN di  USE SIGNAL ; DIRECTION OUTPUT ;
        PORT
        LAYER Metal1 ;
        RECT  87.15 -0.40 87.75 0.30 ;
        END
    END di
    PIN vdd!
        USE power ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        LAYER Metal3 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        END
    END vdd!
    PIN vss!
        USE ground ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        LAYER Metal3 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        END
    END vss!
    OBS
        LAYER Metal1 ;
        RECT  88.35 -0.40 114.75 560.00 ;
        RECT  86.55 0.90 88.35 560.00 ;
        RECT  62.15 -0.40 86.55 560.00 ;
        RECT  60.35 0.90 62.15 560.00 ;
        RECT  27.15 -0.40 60.35 560.00 ;
        RECT  25.35 0.90 27.15 560.00 ;
        RECT  0.25 -0.40 25.35 560.00 ;
        LAYER Metal2 ;
        RECT  0.33 0.33 114.68 559.92 ;
        LAYER Metal3 ;
        RECT  114.65 0.33 114.68 559.92 ;
        RECT  103.70 2.20 114.65 559.92 ;
        RECT  4.05 2.20 14.70 559.92 ;
        RECT  2.20 0.33 4.05 559.92 ;
        RECT  0.33 0.33 2.20 59.75 ;
        RECT  0.33 108.90 2.20 109.60 ;
        RECT  0.33 241.90 2.20 242.60 ;
        RECT  0.33 380.90 2.20 559.92 ;
        RECT  14.70 0.33 103.70 559.92 ;
    END
END iobufs3_16pd_8

MACRO iobufs3_16pu_12
    CLASS PAD ;
    FOREIGN iobufs3_16pu_12  0.00 -38.75 N  ;
    ORIGIN 0.00 39.15 ;
    SIZE 115.00 BY 600.00 ;
    SYMMETRY x y r90 ;
    SITE io_site ;
     PIN en USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  60.95 -0.40 61.55 0.30 ;
        END
    END en
    PIN pad USE SIGNAL ; DIRECTION INOUT ;
        PORT
        LAYER Metal3 ;
        RECT  3.00 383.00 112.00 544.25 ;
        END
    END pad
    PIN do USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  25.95 -0.40 26.55 0.30 ;
        END
    END do
    PIN di  USE SIGNAL ; DIRECTION OUTPUT ;
        PORT
        LAYER Metal1 ;
        RECT  87.15 -0.40 87.75 0.30 ;
        END
    END di
    PIN vdd!
        USE power ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        LAYER Metal3 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        END
    END vdd!
    PIN vss!
        USE ground ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        LAYER Metal3 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        END
    END vss!
    OBS
        LAYER Metal1 ;
        RECT  88.35 -0.40 114.75 560.00 ;
        RECT  86.55 0.90 88.35 560.00 ;
        RECT  62.15 -0.40 86.55 560.00 ;
        RECT  60.35 0.90 62.15 560.00 ;
        RECT  27.15 -0.40 60.35 560.00 ;
        RECT  25.35 0.90 27.15 560.00 ;
        RECT  0.25 -0.40 25.35 560.00 ;
        LAYER Metal2 ;
        RECT  0.33 0.33 114.68 559.92 ;
        LAYER Metal3 ;
        RECT  114.65 0.33 114.68 559.92 ;
        RECT  103.70 2.20 114.65 559.92 ;
        RECT  4.05 2.20 14.70 559.92 ;
        RECT  2.20 0.33 4.05 559.92 ;
        RECT  0.33 0.33 2.20 59.75 ;
        RECT  0.33 108.90 2.20 109.60 ;
        RECT  0.33 241.90 2.20 242.60 ;
        RECT  0.33 380.90 2.20 559.92 ;
        RECT  14.70 0.33 103.70 559.92 ;
    END
END iobufs3_16pu_12

MACRO iobufs3_16pu_4
    CLASS PAD ;
    FOREIGN iobufs3_16pu_4  0.00 -38.75 N  ;
    ORIGIN 0.00 39.15 ;
    SIZE 115.00 BY 600.00 ;
    SYMMETRY x y r90 ;
    SITE io_site ;
     PIN en USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  60.95 -0.40 61.55 0.30 ;
        END
    END en
    PIN pad USE SIGNAL ; DIRECTION INOUT ;
        PORT
        LAYER Metal3 ;
        RECT  3.00 383.00 112.00 544.25 ;
        END
    END pad
    PIN do USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  25.95 -0.40 26.55 0.30 ;
        END
    END do
    PIN di  USE SIGNAL ; DIRECTION OUTPUT ;
        PORT
        LAYER Metal1 ;
        RECT  87.15 -0.40 87.75 0.30 ;
        END
    END di
    PIN vdd!
        USE power ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        LAYER Metal3 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        END
    END vdd!
    PIN vss!
        USE ground ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        LAYER Metal3 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        END
    END vss!
    OBS
        LAYER Metal1 ;
        RECT  88.35 -0.40 114.75 560.00 ;
        RECT  86.55 0.90 88.35 560.00 ;
        RECT  62.15 -0.40 86.55 560.00 ;
        RECT  60.35 0.90 62.15 560.00 ;
        RECT  27.15 -0.40 60.35 560.00 ;
        RECT  25.35 0.90 27.15 560.00 ;
        RECT  0.25 -0.40 25.35 560.00 ;
        LAYER Metal2 ;
        RECT  0.33 0.33 114.68 559.92 ;
        LAYER Metal3 ;
        RECT  114.65 0.33 114.68 559.92 ;
        RECT  103.70 2.20 114.65 559.92 ;
        RECT  4.05 2.20 14.70 559.92 ;
        RECT  2.20 0.33 4.05 559.92 ;
        RECT  0.33 0.33 2.20 59.75 ;
        RECT  0.33 108.90 2.20 109.60 ;
        RECT  0.33 241.90 2.20 242.60 ;
        RECT  0.33 380.90 2.20 559.92 ;
        RECT  14.70 0.33 103.70 559.92 ;
    END
END iobufs3_16pu_4

MACRO iobufs3_16pu_8
    CLASS PAD ;
    FOREIGN iobufs3_16pu_8  0.00 -38.75 N  ;
    ORIGIN 0.00 39.15 ;
    SIZE 115.00 BY 600.00 ;
    SYMMETRY x y r90 ;
    SITE io_site ;
     PIN en USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  60.95 -0.40 61.55 0.30 ;
        END
    END en
    PIN pad USE SIGNAL ; DIRECTION INOUT ;
        PORT
        LAYER Metal3 ;
        RECT  3.00 383.00 112.00 544.25 ;
        END
    END pad
    PIN do USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  25.95 -0.40 26.55 0.30 ;
        END
    END do
    PIN di  USE SIGNAL ; DIRECTION OUTPUT ;
        PORT
        LAYER Metal1 ;
        RECT  87.15 -0.40 87.75 0.30 ;
        END
    END di
    PIN vdd!
        USE power ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        LAYER Metal3 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        END
    END vdd!
    PIN vss!
        USE ground ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        LAYER Metal3 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        END
    END vss!
    OBS
        LAYER Metal1 ;
        RECT  88.35 -0.40 114.75 560.00 ;
        RECT  86.55 0.90 88.35 560.00 ;
        RECT  62.15 -0.40 86.55 560.00 ;
        RECT  60.35 0.90 62.15 560.00 ;
        RECT  27.15 -0.40 60.35 560.00 ;
        RECT  25.35 0.90 27.15 560.00 ;
        RECT  0.25 -0.40 25.35 560.00 ;
        LAYER Metal2 ;
        RECT  0.33 0.33 114.68 559.92 ;
        LAYER Metal3 ;
        RECT  114.65 0.33 114.68 559.92 ;
        RECT  103.70 2.20 114.65 559.92 ;
        RECT  4.05 2.20 14.70 559.92 ;
        RECT  2.20 0.33 4.05 559.92 ;
        RECT  0.33 0.33 2.20 59.75 ;
        RECT  0.33 108.90 2.20 109.60 ;
        RECT  0.33 241.90 2.20 242.60 ;
        RECT  0.33 380.90 2.20 559.92 ;
        RECT  14.70 0.33 103.70 559.92 ;
    END
END iobufs3_16pu_8

MACRO iobufsdv_16_12
    CLASS PAD ;
    FOREIGN iobufsdv_16_12  0.00 -38.75 N  ;
    ORIGIN 0.00 39.15 ;
    SIZE 115.00 BY 600.00 ;
    SYMMETRY x y r90 ;
    SITE io_site ;
     PIN en USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  60.95 -0.40 61.55 0.30 ;
        END
    END en
    PIN pad USE SIGNAL ; DIRECTION INOUT ;
        PORT
        LAYER Metal3 ;
        RECT  3.00 383.00 112.00 544.25 ;
        END
    END pad
    PIN do USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  25.95 -0.40 26.55 0.30 ;
        END
    END do
    PIN di  USE SIGNAL ; DIRECTION OUTPUT ;
        PORT
        LAYER Metal1 ;
        RECT  87.15 -0.40 87.75 0.30 ;
        END
    END di
    PIN vdd!
        USE power ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        LAYER Metal3 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        END
    END vdd!
    PIN vss!
        USE ground ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        LAYER Metal3 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        END
    END vss!
    OBS
        LAYER Metal1 ;
        RECT  88.35 -0.40 114.75 560.00 ;
        RECT  86.55 0.90 88.35 560.00 ;
        RECT  62.15 -0.40 86.55 560.00 ;
        RECT  60.35 0.90 62.15 560.00 ;
        RECT  27.15 -0.40 60.35 560.00 ;
        RECT  25.35 0.90 27.15 560.00 ;
        RECT  0.25 -0.40 25.35 560.00 ;
        LAYER Metal2 ;
        RECT  0.33 0.33 114.68 559.92 ;
        LAYER Metal3 ;
        RECT  114.65 0.33 114.68 559.92 ;
        RECT  103.70 2.20 114.65 559.92 ;
        RECT  4.05 2.20 14.70 559.92 ;
        RECT  2.20 0.33 4.05 559.92 ;
        RECT  0.33 0.33 2.20 59.75 ;
        RECT  0.33 108.90 2.20 109.60 ;
        RECT  0.33 241.90 2.20 242.60 ;
        RECT  0.33 380.90 2.20 559.92 ;
        RECT  14.70 0.33 103.70 559.92 ;
    END
END iobufsdv_16_12

MACRO iobufsdv_16_4
    CLASS PAD ;
    FOREIGN iobufsdv_16_4  0.00 -38.75 N  ;
    ORIGIN 0.00 39.15 ;
    SIZE 115.00 BY 600.00 ;
    SYMMETRY x y r90 ;
    SITE io_site ;
     PIN en USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  60.95 -0.40 61.55 0.30 ;
        END
    END en
    PIN pad USE SIGNAL ; DIRECTION INOUT ;
        PORT
        LAYER Metal3 ;
        RECT  3.00 383.00 112.00 544.25 ;
        END
    END pad
    PIN do USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  25.95 -0.40 26.55 0.30 ;
        END
    END do
    PIN di  USE SIGNAL ; DIRECTION OUTPUT ;
        PORT
        LAYER Metal1 ;
        RECT  87.15 -0.40 87.75 0.30 ;
        END
    END di
    PIN vdd!
        USE power ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        LAYER Metal3 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        END
    END vdd!
    PIN vss!
        USE ground ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        LAYER Metal3 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        END
    END vss!
    OBS
        LAYER Metal1 ;
        RECT  88.35 -0.40 114.75 560.00 ;
        RECT  86.55 0.90 88.35 560.00 ;
        RECT  62.15 -0.40 86.55 560.00 ;
        RECT  60.35 0.90 62.15 560.00 ;
        RECT  27.15 -0.40 60.35 560.00 ;
        RECT  25.35 0.90 27.15 560.00 ;
        RECT  0.25 -0.40 25.35 560.00 ;
        LAYER Metal2 ;
        RECT  0.33 0.33 114.68 559.92 ;
        LAYER Metal3 ;
        RECT  114.65 0.33 114.68 559.92 ;
        RECT  103.70 2.20 114.65 559.92 ;
        RECT  4.05 2.20 14.70 559.92 ;
        RECT  2.20 0.33 4.05 559.92 ;
        RECT  0.33 0.33 2.20 59.75 ;
        RECT  0.33 108.90 2.20 109.60 ;
        RECT  0.33 241.90 2.20 242.60 ;
        RECT  0.33 380.90 2.20 559.92 ;
        RECT  14.70 0.33 103.70 559.92 ;
    END
END iobufsdv_16_4

MACRO iobufsdv_16_8
    CLASS PAD ;
    FOREIGN iobufsdv_16_8  0.00 -38.75 N  ;
    ORIGIN 0.00 39.15 ;
    SIZE 115.00 BY 600.00 ;
    SYMMETRY x y r90 ;
    SITE io_site ;
     PIN en USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  60.95 -0.40 61.55 0.30 ;
        END
    END en
    PIN pad USE SIGNAL ; DIRECTION INOUT ;
        PORT
        LAYER Metal3 ;
        RECT  3.00 383.00 112.00 544.25 ;
        END
    END pad
    PIN do USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  25.95 -0.40 26.55 0.30 ;
        END
    END do
    PIN di  USE SIGNAL ; DIRECTION OUTPUT ;
        PORT
        LAYER Metal1 ;
        RECT  87.15 -0.40 87.75 0.30 ;
        END
    END di
    PIN vdd!
        USE power ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        LAYER Metal3 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        END
    END vdd!
    PIN vss!
        USE ground ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        LAYER Metal3 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        END
    END vss!
    OBS
        LAYER Metal1 ;
        RECT  88.35 -0.40 114.75 560.00 ;
        RECT  86.55 0.90 88.35 560.00 ;
        RECT  62.15 -0.40 86.55 560.00 ;
        RECT  60.35 0.90 62.15 560.00 ;
        RECT  27.15 -0.40 60.35 560.00 ;
        RECT  25.35 0.90 27.15 560.00 ;
        RECT  0.25 -0.40 25.35 560.00 ;
        LAYER Metal2 ;
        RECT  0.33 0.33 114.68 559.92 ;
        LAYER Metal3 ;
        RECT  114.65 0.33 114.68 559.92 ;
        RECT  103.70 2.20 114.65 559.92 ;
        RECT  4.05 2.20 14.70 559.92 ;
        RECT  2.20 0.33 4.05 559.92 ;
        RECT  0.33 0.33 2.20 59.75 ;
        RECT  0.33 108.90 2.20 109.60 ;
        RECT  0.33 241.90 2.20 242.60 ;
        RECT  0.33 380.90 2.20 559.92 ;
        RECT  14.70 0.33 103.70 559.92 ;
    END
END iobufsdv_16_8

MACRO iobufsdv_16pd_12
    CLASS PAD ;
    FOREIGN iobufsdv_16pd_12  0.00 -38.75 N  ;
    ORIGIN 0.00 39.15 ;
    SIZE 115.00 BY 600.00 ;
    SYMMETRY x y r90 ;
    SITE io_site ;
     PIN en USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  60.95 -0.40 61.55 0.30 ;
        END
    END en
    PIN pad USE SIGNAL ; DIRECTION INOUT ;
        PORT
        LAYER Metal3 ;
        RECT  3.00 383.00 112.00 544.25 ;
        END
    END pad
    PIN do USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  25.95 -0.40 26.55 0.30 ;
        END
    END do
    PIN di  USE SIGNAL ; DIRECTION OUTPUT ;
        PORT
        LAYER Metal1 ;
        RECT  87.15 -0.40 87.75 0.30 ;
        END
    END di
    PIN vdd!
        USE power ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        LAYER Metal3 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        END
    END vdd!
    PIN vss!
        USE ground ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        LAYER Metal3 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        END
    END vss!
    OBS
        LAYER Metal1 ;
        RECT  88.35 -0.40 114.75 560.00 ;
        RECT  86.55 0.90 88.35 560.00 ;
        RECT  62.15 -0.40 86.55 560.00 ;
        RECT  60.35 0.90 62.15 560.00 ;
        RECT  27.15 -0.40 60.35 560.00 ;
        RECT  25.35 0.90 27.15 560.00 ;
        RECT  0.25 -0.40 25.35 560.00 ;
        LAYER Metal2 ;
        RECT  0.33 0.33 114.68 559.92 ;
        LAYER Metal3 ;
        RECT  114.65 0.33 114.68 559.92 ;
        RECT  103.70 2.20 114.65 559.92 ;
        RECT  4.05 2.20 14.70 559.92 ;
        RECT  2.20 0.33 4.05 559.92 ;
        RECT  0.33 0.33 2.20 59.75 ;
        RECT  0.33 108.90 2.20 109.60 ;
        RECT  0.33 241.90 2.20 242.60 ;
        RECT  0.33 380.90 2.20 559.92 ;
        RECT  14.70 0.33 103.70 559.92 ;
    END
END iobufsdv_16pd_12

MACRO iobufsdv_16pd_4
    CLASS PAD ;
    FOREIGN iobufsdv_16pd_4  0.00 -38.75 N  ;
    ORIGIN 0.00 39.15 ;
    SIZE 115.00 BY 600.00 ;
    SYMMETRY x y r90 ;
    SITE io_site ;
     PIN en USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  60.95 -0.40 61.55 0.30 ;
        END
    END en
    PIN pad USE SIGNAL ; DIRECTION INOUT ;
        PORT
        LAYER Metal3 ;
        RECT  3.00 383.00 112.00 544.25 ;
        END
    END pad
    PIN do USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  25.95 -0.40 26.55 0.30 ;
        END
    END do
    PIN di  USE SIGNAL ; DIRECTION OUTPUT ;
        PORT
        LAYER Metal1 ;
        RECT  87.15 -0.40 87.75 0.30 ;
        END
    END di
    PIN vdd!
        USE power ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        LAYER Metal3 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        END
    END vdd!
    PIN vss!
        USE ground ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        LAYER Metal3 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        END
    END vss!
    OBS
        LAYER Metal1 ;
        RECT  88.35 -0.40 114.75 560.00 ;
        RECT  86.55 0.90 88.35 560.00 ;
        RECT  62.15 -0.40 86.55 560.00 ;
        RECT  60.35 0.90 62.15 560.00 ;
        RECT  27.15 -0.40 60.35 560.00 ;
        RECT  25.35 0.90 27.15 560.00 ;
        RECT  0.25 -0.40 25.35 560.00 ;
        LAYER Metal2 ;
        RECT  0.33 0.33 114.68 559.92 ;
        LAYER Metal3 ;
        RECT  114.65 0.33 114.68 559.92 ;
        RECT  103.70 2.20 114.65 559.92 ;
        RECT  4.05 2.20 14.70 559.92 ;
        RECT  2.20 0.33 4.05 559.92 ;
        RECT  0.33 0.33 2.20 59.75 ;
        RECT  0.33 108.90 2.20 109.60 ;
        RECT  0.33 241.90 2.20 242.60 ;
        RECT  0.33 380.90 2.20 559.92 ;
        RECT  14.70 0.33 103.70 559.92 ;
    END
END iobufsdv_16pd_4

MACRO iobufsdv_16pd_8
    CLASS PAD ;
    FOREIGN iobufsdv_16pd_8  0.00 -38.75 N  ;
    ORIGIN 0.00 39.15 ;
    SIZE 115.00 BY 600.00 ;
    SYMMETRY x y r90 ;
    SITE io_site ;
     PIN en USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  60.95 -0.40 61.55 0.30 ;
        END
    END en
    PIN pad USE SIGNAL ; DIRECTION INOUT ;
        PORT
        LAYER Metal3 ;
        RECT  3.00 383.00 112.00 544.25 ;
        END
    END pad
    PIN do USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  25.95 -0.40 26.55 0.30 ;
        END
    END do
    PIN di  USE SIGNAL ; DIRECTION OUTPUT ;
        PORT
        LAYER Metal1 ;
        RECT  87.15 -0.40 87.75 0.30 ;
        END
    END di
    PIN vdd!
        USE power ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        LAYER Metal3 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        END
    END vdd!
    PIN vss!
        USE ground ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        LAYER Metal3 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        END
    END vss!
    OBS
        LAYER Metal1 ;
        RECT  88.35 -0.40 114.75 560.00 ;
        RECT  86.55 0.90 88.35 560.00 ;
        RECT  62.15 -0.40 86.55 560.00 ;
        RECT  60.35 0.90 62.15 560.00 ;
        RECT  27.15 -0.40 60.35 560.00 ;
        RECT  25.35 0.90 27.15 560.00 ;
        RECT  0.25 -0.40 25.35 560.00 ;
        LAYER Metal2 ;
        RECT  0.33 0.33 114.68 559.92 ;
        LAYER Metal3 ;
        RECT  114.65 0.33 114.68 559.92 ;
        RECT  103.70 2.20 114.65 559.92 ;
        RECT  4.05 2.20 14.70 559.92 ;
        RECT  2.20 0.33 4.05 559.92 ;
        RECT  0.33 0.33 2.20 59.75 ;
        RECT  0.33 108.90 2.20 109.60 ;
        RECT  0.33 241.90 2.20 242.60 ;
        RECT  0.33 380.90 2.20 559.92 ;
        RECT  14.70 0.33 103.70 559.92 ;
    END
END iobufsdv_16pd_8

MACRO iobufsdv_16pu_12
    CLASS PAD ;
    FOREIGN iobufsdv_16pu_12  0.00 -38.75 N  ;
    ORIGIN 0.00 39.15 ;
    SIZE 115.00 BY 600.00 ;
    SYMMETRY x y r90 ;
    SITE io_site ;
     PIN en USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  60.95 -0.40 61.55 0.30 ;
        END
    END en
    PIN pad USE SIGNAL ; DIRECTION INOUT ;
        PORT
        LAYER Metal3 ;
        RECT  3.00 383.00 112.00 544.25 ;
        END
    END pad
    PIN do USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  25.95 -0.40 26.55 0.30 ;
        END
    END do
    PIN di  USE SIGNAL ; DIRECTION OUTPUT ;
        PORT
        LAYER Metal1 ;
        RECT  87.15 -0.40 87.75 0.30 ;
        END
    END di
    PIN vdd!
        USE power ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        LAYER Metal3 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        END
    END vdd!
    PIN vss!
        USE ground ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        LAYER Metal3 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        END
    END vss!
    OBS
        LAYER Metal1 ;
        RECT  88.35 -0.40 114.75 560.00 ;
        RECT  86.55 0.90 88.35 560.00 ;
        RECT  62.15 -0.40 86.55 560.00 ;
        RECT  60.35 0.90 62.15 560.00 ;
        RECT  27.15 -0.40 60.35 560.00 ;
        RECT  25.35 0.90 27.15 560.00 ;
        RECT  0.25 -0.40 25.35 560.00 ;
        LAYER Metal2 ;
        RECT  0.33 0.33 114.68 559.92 ;
        LAYER Metal3 ;
        RECT  114.65 0.33 114.68 559.92 ;
        RECT  103.70 2.20 114.65 559.92 ;
        RECT  4.05 2.20 14.70 559.92 ;
        RECT  2.20 0.33 4.05 559.92 ;
        RECT  0.33 0.33 2.20 59.75 ;
        RECT  0.33 108.90 2.20 109.60 ;
        RECT  0.33 241.90 2.20 242.60 ;
        RECT  0.33 380.90 2.20 559.92 ;
        RECT  14.70 0.33 103.70 559.92 ;
    END
END iobufsdv_16pu_12

MACRO iobufsdv_16pu_4
    CLASS PAD ;
    FOREIGN iobufsdv_16pu_4  0.00 -38.75 N  ;
    ORIGIN 0.00 39.15 ;
    SIZE 115.00 BY 600.00 ;
    SYMMETRY x y r90 ;
    SITE io_site ;
     PIN en USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  60.95 -0.40 61.55 0.30 ;
        END
    END en
    PIN pad USE SIGNAL ; DIRECTION INOUT ;
        PORT
        LAYER Metal3 ;
        RECT  3.00 383.00 112.00 544.25 ;
        END
    END pad
    PIN do USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  25.95 -0.40 26.55 0.30 ;
        END
    END do
    PIN di  USE SIGNAL ; DIRECTION OUTPUT ;
        PORT
        LAYER Metal1 ;
        RECT  87.15 -0.40 87.75 0.30 ;
        END
    END di
    PIN vdd!
        USE power ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        LAYER Metal3 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        END
    END vdd!
    PIN vss!
        USE ground ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        LAYER Metal3 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        END
    END vss!
    OBS
        LAYER Metal1 ;
        RECT  88.35 -0.40 114.75 560.00 ;
        RECT  86.55 0.90 88.35 560.00 ;
        RECT  62.15 -0.40 86.55 560.00 ;
        RECT  60.35 0.90 62.15 560.00 ;
        RECT  27.15 -0.40 60.35 560.00 ;
        RECT  25.35 0.90 27.15 560.00 ;
        RECT  0.25 -0.40 25.35 560.00 ;
        LAYER Metal2 ;
        RECT  0.33 0.33 114.68 559.92 ;
        LAYER Metal3 ;
        RECT  114.65 0.33 114.68 559.92 ;
        RECT  103.70 2.20 114.65 559.92 ;
        RECT  4.05 2.20 14.70 559.92 ;
        RECT  2.20 0.33 4.05 559.92 ;
        RECT  0.33 0.33 2.20 59.75 ;
        RECT  0.33 108.90 2.20 109.60 ;
        RECT  0.33 241.90 2.20 242.60 ;
        RECT  0.33 380.90 2.20 559.92 ;
        RECT  14.70 0.33 103.70 559.92 ;
    END
END iobufsdv_16pu_4

MACRO iobufsdv_16pu_8
    CLASS PAD ;
    FOREIGN iobufsdv_16pu_8  0.00 -38.75 N  ;
    ORIGIN 0.00 39.15 ;
    SIZE 115.00 BY 600.00 ;
    SYMMETRY x y r90 ;
    SITE io_site ;
     PIN en USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  60.95 -0.40 61.55 0.30 ;
        END
    END en
    PIN pad USE SIGNAL ; DIRECTION INOUT ;
        PORT
        LAYER Metal3 ;
        RECT  3.00 383.00 112.00 544.25 ;
        END
    END pad
    PIN do USE SIGNAL ; DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  25.95 -0.40 26.55 0.30 ;
        END
    END do
    PIN di  USE SIGNAL ; DIRECTION OUTPUT ;
        PORT
        LAYER Metal1 ;
        RECT  87.15 -0.40 87.75 0.30 ;
        END
    END di
    PIN vdd!
        USE power ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        LAYER Metal3 ;
        RECT  104.35 -0.40 114.00 1.55 ;
        END
    END vdd!
    PIN vss!
        USE ground ;  DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        LAYER Metal3 ;
         RECT  4.75 -0.40 14.05 1.55 ;
        END
    END vss!
    OBS
        LAYER Metal1 ;
        RECT  88.35 -0.40 114.75 560.00 ;
        RECT  86.55 0.90 88.35 560.00 ;
        RECT  62.15 -0.40 86.55 560.00 ;
        RECT  60.35 0.90 62.15 560.00 ;
        RECT  27.15 -0.40 60.35 560.00 ;
        RECT  25.35 0.90 27.15 560.00 ;
        RECT  0.25 -0.40 25.35 560.00 ;
        LAYER Metal2 ;
        RECT  0.33 0.33 114.68 559.92 ;
        LAYER Metal3 ;
        RECT  114.65 0.33 114.68 559.92 ;
        RECT  103.70 2.20 114.65 559.92 ;
        RECT  4.05 2.20 14.70 559.92 ;
        RECT  2.20 0.33 4.05 559.92 ;
        RECT  0.33 0.33 2.20 59.75 ;
        RECT  0.33 108.90 2.20 109.60 ;
        RECT  0.33 241.90 2.20 242.60 ;
        RECT  0.33 380.90 2.20 559.92 ;
        RECT  14.70 0.33 103.70 559.92 ;
    END
END iobufsdv_16pu_8

MACRO llcnr_sep
    CLASS ENDCAP BOTTOMLEFT ;
    FOREIGN llcnr_sep 0.00 0.00  ;
    ORIGIN 0.00  0.00 ;
    SIZE 600.00 BY 600.00 ;
    SYMMETRY x y r90 ;
    SITE io_corner ;
    OBS
        LAYER Metal1 ;
        RECT  0.25 0.25 598.75 598.75 ;
        LAYER Metal2 ;
        RECT  0.33 0.33 598.67 598.67 ;
        LAYER Metal3 ;
        RECT  0.33 0.33 598.67 598.67 ;
        LAYER Metal4 ;
        RECT  0.33 0.33 598.67 598.67 ;
        LAYER Metal5 ;
        RECT  0.33 0.33 598.67 598.67 ;
    END
END llcnr_sep

MACRO llcnr_tie
    CLASS ENDCAP BOTTOMLEFT ;
    FOREIGN llcnr_tie 0.00 0.00  ;
    ORIGIN 0.00  0.00 ;
    SIZE 600.00 BY 600.00 ;
    SYMMETRY x y r90 ;
    SITE io_corner ;
    OBS
        LAYER Metal1 ;
        RECT  0.25 0.25 598.75 598.75 ;
        LAYER Metal2 ;
        RECT  0.33 0.33 598.67 598.67 ;
        LAYER Metal3 ;
        RECT  0.33 0.33 598.67 598.67 ;
        LAYER Metal4 ;
        RECT  0.33 0.33 598.67 598.67 ;
        LAYER Metal5 ;
        RECT  0.33 0.33 598.67 598.67 ;
    END
END llcnr_tie

MACRO lrcnr_sep
    CLASS ENDCAP BOTTOMLEFT ;
    FOREIGN lrcnr_sep 0.00 0.00  ;
    ORIGIN 0.00  0.00 ;
    SIZE 600.00 BY 600.00 ;
    SYMMETRY x y r90 ;
    SITE io_corner ;
    OBS
        LAYER Metal1 ;
        RECT  0.25 0.25 598.75 598.75 ;
        LAYER Metal2 ;
        RECT  0.33 0.33 598.67 598.67 ;
        LAYER Metal3 ;
        RECT  0.33 0.33 598.67 598.67 ;
        LAYER Metal4 ;
        RECT  0.33 0.33 598.67 598.67 ;
        LAYER Metal5 ;
        RECT  0.33 0.33 598.67 598.67 ;
    END
END lrcnr_sep

MACRO lrcnr_tie
    CLASS ENDCAP BOTTOMLEFT ;
    FOREIGN lrcnr_tie 0.00 0.00  ;
    ORIGIN 0.00  0.00 ;
    SIZE 600.00 BY 600.00 ;
    SYMMETRY x y r90 ;
    SITE io_corner ;
    OBS
        LAYER Metal1 ;
        RECT  0.25 0.25 598.75 598.75 ;
        LAYER Metal2 ;
        RECT  0.33 0.33 598.67 598.67 ;
        LAYER Metal3 ;
        RECT  0.33 0.33 598.67 598.67 ;
        LAYER Metal4 ;
        RECT  0.33 0.33 598.67 598.67 ;
        LAYER Metal5 ;
        RECT  0.33 0.33 598.67 598.67 ;
    END
END lrcnr_tie

MACRO outvdd
    CLASS PAD ;
    FOREIGN outvdd  0.00 -38.75 N  ;
    ORIGIN 0.00  39.15 ;
    SIZE 115.00 BY 600.00 ;
    SYMMETRY x y r90 ;
    SITE io_site ;
    PIN pad USE POWER ; DIRECTION INPUT ;
        PORT
        LAYER Metal5 ;
        RECT  3.00 383.00 112.00 544.25 ;
        END
    END pad
    OBS
        LAYER Metal1 ;
        RECT  0.25 -0.40 114.75 560.00 ;
        LAYER Metal2 ;
        RECT  0.33 0.33 114.68 559.92 ;
        LAYER Metal3 ;
        RECT  0.33 0.33 114.68 559.92 ;
        LAYER Metal4 ;
        RECT  0.33 0.33 114.68 559.92 ;
        LAYER Metal5 ;
        RECT  0.33 0.33 114.68 559.92 ;
    END
END outvdd

MACRO outvss
    CLASS PAD ;
    FOREIGN outvss  0.00 -38.75 N  ;
    ORIGIN 0.00 39.15 ;
    SIZE 115.00 BY 600.00 ;
    SYMMETRY x y r90 ;
    SITE io_site ;
    PIN pad USE power ; DIRECTION INPUT ;
        PORT
        LAYER Metal5 ;
        RECT  3.00 383.00 112.00 544.25 ;
        END
    END pad
    OBS
        LAYER Metal1 ;
        RECT  0.25 -0.40 114.75 560.00 ;
        LAYER Metal2 ;
        RECT  0.33 0.33 114.68 559.92 ;
        LAYER Metal3 ;
        RECT  0.33 0.33 114.68 559.92 ;
        LAYER Metal4 ;
        RECT  0.33 0.33 114.68 559.92 ;
        LAYER Metal5 ;
        RECT  0.33 0.33 114.68 559.92 ;
    END
END outvss

MACRO ulcnr_sep
    CLASS ENDCAP BOTTOMLEFT ;
    FOREIGN ulcnr_sep 0.00 0.00  ;
    ORIGIN 0.00  0.00 ;
    SIZE 600.00 BY 600.00 ;
    SYMMETRY x y r90 ;
    SITE io_corner ;
    OBS
        LAYER Metal1 ;
        RECT  0.25 0.25 598.75 598.75 ;
        LAYER Metal2 ;
        RECT  0.33 0.33 598.67 598.67 ;
        LAYER Metal3 ;
        RECT  0.33 0.33 598.67 598.67 ;
        LAYER Metal4 ;
        RECT  0.33 0.33 598.67 598.67 ;
        LAYER Metal5 ;
        RECT  0.33 0.33 598.67 598.67 ;
    END
END ulcnr_sep

MACRO ulcnr_tie
    CLASS ENDCAP BOTTOMLEFT ;
    FOREIGN ulcnr_tie 0.00 0.00  ;
    ORIGIN 0.00  0.00 ;
    SIZE 600.00 BY 600.00 ;
    SYMMETRY x y r90 ;
    SITE io_corner ;
    OBS
        LAYER Metal1 ;
        RECT  0.25 0.25 598.75 598.75 ;
        LAYER Metal2 ;
        RECT  0.33 0.33 598.67 598.67 ;
        LAYER Metal3 ;
        RECT  0.33 0.33 598.67 598.67 ;
        LAYER Metal4 ;
        RECT  0.33 0.33 598.67 598.67 ;
        LAYER Metal5 ;
        RECT  0.33 0.33 598.67 598.67 ;
    END
END ulcnr_tie

MACRO urcnr_sep
    CLASS ENDCAP BOTTOMLEFT ;
    FOREIGN urcnr_sep 0.00 0.00  ;
    ORIGIN 0.00  0.00 ;
    SIZE 600.00 BY 600.00 ;
    SYMMETRY x y r90 ;
    SITE io_corner ;
    OBS
        LAYER Metal1 ;
        RECT  0.25 0.25 598.75 598.75 ;
        LAYER Metal2 ;
        RECT  0.33 0.33 598.67 598.67 ;
        LAYER Metal3 ;
        RECT  0.33 0.33 598.67 598.67 ;
        LAYER Metal4 ;
        RECT  0.33 0.33 598.67 598.67 ;
        LAYER Metal5 ;
        RECT  0.33 0.33 598.67 598.67 ;
    END
END urcnr_sep

MACRO urcnr_tie
    CLASS ENDCAP BOTTOMLEFT ;
    FOREIGN urcnr_tie 0.00 0.00  ;
    ORIGIN 0.00  0.00 ;
    SIZE 600.00 BY 600.00 ;
    SYMMETRY x y r90 ;
    SITE io_corner ;
    OBS
        LAYER Metal1 ;
        RECT  0.25 0.25 598.75 598.75 ;
        LAYER Metal2 ;
        RECT  0.33 0.33 598.67 598.67 ;
        LAYER Metal3 ;
        RECT  0.33 0.33 598.67 598.67 ;
        LAYER Metal4 ;
        RECT  0.33 0.33 598.67 598.67 ;
        LAYER Metal5 ;
        RECT  0.33 0.33 598.67 598.67 ;
    END
END urcnr_tie

#END LIBRARY
#7.3.03 u.j. + g.p. from GDS to lef
# correction 13.11.03 u.j.

#VERSION 5.4 ;

MACRO sram2k_pin
    CLASS BLOCK ;
    FOREIGN sram2k_pin 0 0 N ;
    SYMMETRY X Y r90 ;
    SIZE  1682.40 BY 949.55 ;
    SITE core ;
    PIN vdd!
        USE power ;  
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  1676.4 34.4 1682.4 65.65 ; 
        RECT  1676.4 75.5  1682.4 81.75 ;
        RECT  1676.4 867.5  1682.4 873.75 ;
        RECT  1676.4 883.75  1682.4 915.0 ;
        RECT  0.0 883.75  6.0 915.0 ;
        RECT  0.0 867.5  6.0 873.75 ;
        RECT  0.0 774.0  6.0 780.25 ;
        RECT  0.0 75.5  6.0 81.75 ; 
        RECT  0.0 34.4  6.0 65.65 ;
        END
    END vdd! 
    PIN vss!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ; 
        RECT 1676.4 916.25 1682.4 947.5 ;
        RECT 1676.4 875.0 1682.4 881.25 ;
        RECT 1676.4 68.0 1682.4 74.25 ;
        RECT 1676.4 1.55 1682.4 32.8 ;
        RECT 0.0 1.55 6.0 32.8 ;
        RECT 0.0 68.0 6.0 74.25 ;
        RECT 0.0 781.5 6.0 787.75 ;
        RECT 0.0 875.0 6.0 881.25 ;
        RECT 0.0 916.25 6.0 947.5 ; 
        END
    END vss! 

PIN oen3
	DIRECTION INPUT ;
	PORT
	LAYER Metal3 ;
	RECT 1328.15 948.55 1330.15 949.55 ;
	END
END oen3

PIN oen2
	DIRECTION INPUT ;
	PORT
	LAYER Metal3 ;
	RECT 980.55 948.55 982.55 949.55 ;
	END
END oen2

PIN oen1
	DIRECTION INPUT ;
	PORT
	LAYER Metal3 ;
	RECT 632.95 948.55 634.95 949.55 ;
	END
END oen1

PIN oen0
	DIRECTION INPUT ;
	PORT
	LAYER Metal3 ;
	RECT 285.35 948.55 287.35 949.55 ;
	END
END oen0

PIN iwen3
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 1126.25 0.0 1128.25 0.6 ;
	END
END iwen3

PIN iwen2
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 1119.75 0.0 1121.75 0.6 ;
	END
END iwen2

PIN iwen1
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 1088.55 0.0 1090.55 0.6 ;
	END
END iwen1

PIN iwen0
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 1080.75 0.0 1082.75 0.6 ;
	END
END iwen0

PIN di31
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 1039.15 0.0 1041.15 0.6 ;
	END
END di31

PIN di30
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 1032.65 0.0 1034.65 0.6 ;
	END
END di30

PIN di29
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 1001.45 0.0 1003.45 0.6 ;
	END
END di29

PIN di28
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 993.65 0.0 995.65 0.6 ;
	END
END di28

PIN di27
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 952.05 0.0 954.05 0.6 ;
	END
END di27

PIN di26
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 945.55 0.0 947.55 0.6 ;
	END
END di26

PIN di25
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 914.35 0.0 916.35 0.6 ;
	END
END di25

PIN di24
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 907.85 0.0 909.85 0.6 ;
	END
END di24

PIN di23
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 866.25 0.0 868.25 0.6 ;
	END
END di23

PIN di22
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 858.45 0.0 860.45 0.6 ;
	END
END di22

PIN di21
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 827.25 0.0 829.25 0.6 ;
	END
END di21

PIN di20
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 820.75 0.0 822.75 0.6 ;
	END
END di20

PIN di19
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 779.15 0.0 781.15 0.6 ;
	END
END di19

PIN di18
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 771.35 0.0 773.35 0.6 ;
	END
END di18

PIN di17
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 740.15 0.0 742.15 0.6 ;
	END
END di17

PIN di16
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 733.65 0.0 735.65 0.6 ;
	END
END di16

PIN di15
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 692.05 0.0 694.05 0.6 ;
	END
END di15

PIN di14
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 684.25 0.0 686.25 0.6 ;
	END
END di14

PIN di13
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 654.35 0.0 656.35 0.6 ;
	END
END di13

PIN di12
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 646.55 0.0 648.55 0.6 ;
	END
END di12

PIN di11
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 604.95 0.0 606.95 0.6 ;
	END
END di11

PIN di10
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 597.15 0.0 599.15 0.6 ;
	END
END di10

PIN di9
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 567.25 0.0 569.25 0.6 ;
	END
END di9

PIN di8
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 559.45 0.0 561.45 0.6 ;
	END
END di8

PIN di7
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 517.85 0.0 519.85 0.6 ;
	END
END di7

PIN di6
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 511.35 0.0 513.35 0.6 ;
	END
END di6

PIN di5
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 480.15 0.0 482.15 0.6 ;
	END
END di5

PIN di4
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 472.35 0.0 474.35 0.6 ;
	END
END di4

PIN di3
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 430.75 0.0 432.75 0.6 ;
	END
END di3

PIN di2
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 424.25 0.0 426.25 0.6 ;
	END
END di2

PIN di1
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 393.05 0.0 395.05 0.6 ;
	END
END di1

PIN di0
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 385.25 0.0 387.25 0.6 ;
	END
END di0

PIN a0
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 161.65 0.0 163.65 0.6 ;
	END
END a0

PIN a1
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 144.75 0.0 146.75 0.6 ; 
	END
END a1

PIN a2
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 134.35 0.0 136.35 0.6 ;
	END
END a2


PIN a3
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 93.75 0.0 95.75 0.6 ;
	END
END a3

PIN wrb
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 80.45 0.0 82.45 0.6 ;
	END
END wrb

PIN ceb
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 77.75 0.0 79.75 0.6 ;
	END
END ceb

PIN clk
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 66.75 0.0 68.75 0.6 ;
	END
END clk

PIN a4
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 59.35 0.0 61.35 0.6 ;
	END
END a4

PIN a5
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 55.95 0.0 57.95 0.6 ;
	END
END a5

PIN a6
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 51.15 0.0 53.15 0.6 ;
	END
END a6

PIN a7
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 42.05 0.0 44.05 0.6 ;
	END
END a7

PIN a8
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 36.85 0.0 38.85 0.6 ;
	END
END a8

PIN do0
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 301.55 948.55 303.45 949.55 ;
	END
END do0

PIN do1
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 342.75 948.55 344.65 949.55 ;
	END
END do1

PIN do2
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 388.45 948.55 390.35 949.55 ;
	END
END do2

PIN do3
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 429.65 948.55 431.55 949.55 ;
	END
END do3

PIN do4
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 475.35 948.55 477.25 949.55 ;
	END
END do4

PIN do5
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 516.55 948.55 518.45 949.55 ;
	END
END do5

PIN do6
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 562.25 948.55 564.15 949.55 ;
	END
END do6

PIN do7
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 603.45 948.55 605.35 949.55 ;
	END
END do7

PIN do8
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 649.15 948.55 651.05 949.55 ;
	END
END do8

PIN do9
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 690.35 948.55 692.25 949.55 ;
	END
END do9

PIN do10
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 736.05 948.55 737.95 949.55 ;
	END
END do10

PIN do11
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 777.25 948.55 779.15 949.55 ;
	END
END do11

PIN do12
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 822.95 948.55 824.85 949.55 ;
	END
END do12

PIN do13
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 864.15 948.55 866.05 949.55 ;
	END
END do13

PIN do14
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 909.85 948.55 911.75 949.55 ;
	END
END do14

PIN do15
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 951.05 948.55 952.95 949.55 ;
	END
END do15

PIN do16
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 996.75 948.55 998.65 949.55 ;
	END
END do16

PIN do17
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 1037.95 948.55 1039.85 949.55 ;
	END
END do17

PIN do18
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 1083.65 948.55 1085.55 949.55 ;
	END
END do18

PIN do19
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 1124.85 948.55 1126.75 949.55 ;
	END
END do19

PIN do20
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 1170.55 948.55 1172.45 949.55 ;
	END
END do20

PIN do21
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 1211.75 948.55 1213.65 949.55 ;
	END
END do21

PIN do22
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 1257.45 948.55 1259.35 949.55 ;
	END
END do22

PIN do23
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 1298.65 948.55 1300.55 949.55 ;
	END
END do23

PIN do24
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 1344.35 948.55 1346.25 949.55 ;
	END
END do24

PIN do25
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 1385.55 948.55 1387.45 949.55 ;
	END
END do25

PIN do26
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 1431.25 948.55 1433.15 949.55 ;
	END
END do26

PIN do27
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 1472.45 948.55 1474.35 949.55 ;
	END
END do27

PIN do28
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 1518.15 948.55 1520.05 949.55 ;
	END
END do28

PIN do29
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 1559.35 948.55 1561.25 949.55 ;
	END
END do29

PIN do30
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 1605.05 948.55 1606.95 949.55 ;
	END
END do30

      PIN do31
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 1646.25 948.55 1648.15 949.55 ;
	END
      END do31
      OBS
        LAYER Metal1 ;
	RECT 1.40 1.40 1681.00 948.15 ;
        LAYER Metal2 ;
	RECT 1.40 1.40 1681.00 948.15 ;
        LAYER Metal3 ;
	RECT 1.40 1.40 1681.00 948.15 ;
        LAYER Metal4 ;
	RECT 1.40 1.40 1681.00 948.15 ;
      END
END sram2k_pin

#10.3.03 h.f. + u.j. + g.p. from GDS to lef
# correction 13.11.03 u.j.
#VERSION 5.4 ;

MACRO sram8k_pin
    CLASS BLOCK ;
    FOREIGN sram8k_pin 0 0 N ;
    SYMMETRY X Y r90 ;
    SIZE   1682.558 BY 2130.35 ;
    SITE core ;
    PIN vdd!
        USE power ;  
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT 1676.4 34.4 1682.4 65.65 ;
        RECT 1676.4 75.5 1682.4 81.75 ;
        RECT 1676.4 955.0 1682.4 961.25 ;
        RECT 1676.4 1845.0 1682.4 1851.25 ;
       RECT 1676.4 2048.75 1682.4 2055.0 ;
       RECT 1676.4 2065.0 1682.4 2096.25 ;
       RECT 0.0 2065.0 6.0 2096.25 ;
       RECT 0.0 2048.75 6.0 2055.0 ;
       RECT 0.0 1489.0 6.0 1495.25 ;
       RECT 0.0 774.0 6.0 780.25 ;
       RECT 0.0 75.5 6.0 81.75 ;
       RECT 0.0 34.4 6.0 65.65 ;
       END
    END vdd! 
    PIN vss!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ; 
        RECT 0.0 781.5 6.0 787.75 ;
        RECT 0.0 1496.5 6.0 1502.75 ;
        RECT 0.0 2056.25 6.0 2062.5 ;
        RECT 0.0 68.0 6.0 74.25 ;
        RECT 0.0 1.55 6.0 32.8 ;
        RECT 1676.4 1.55 1682.4 32.8 ;
        RECT 1676.4 68.0 1682.4 74.25 ;
        RECT 1676.4 962.5 1682.4 968.75 ;
        RECT 1676.4 1852.5 1682.4 1858.75 ;
        RECT 1676.4 2056.25 1682.4 2062.5 ;
        RECT 1676.4 2097.5 1682.4 2128.75 ;
        RECT 0.0 2097.5 6.0 2128.75 ;
        END
     END vss!



PIN oen3
	DIRECTION INPUT ;
	PORT
	LAYER Metal3 ;
	RECT 1328.15 2129.1 1330.15 2130.35 ;
	END
END oen3

PIN oen2
	DIRECTION INPUT ;
	PORT
	LAYER Metal3 ;
	RECT 980.55 2129.1 982.55 2130.35 ;
	END
END oen2

PIN oen1
	DIRECTION INPUT ;
	PORT
	LAYER Metal3 ;
	RECT 632.95 2129.1 634.95 2130.35 ;
	END
END oen1

PIN oen0
	DIRECTION INPUT ;
	PORT
	LAYER Metal3 ;
	RECT 285.35 2129.1 287.35 2130.35 ;
	END
END oen0

PIN do31
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 1646.25 2129.1 1648.15 2130.35 ;
	END
END do31

PIN do30
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 1605.05 2129.1 1606.95 2130.35 ;
	END
END do30

PIN do29
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 1559.35 2129.1 1561.25 2130.35 ;
	END
END do29

PIN do28
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 1518.15 2129.1 1520.05 2130.35 ;
	END
END do28

PIN do27
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 1472.45 2129.1 1474.35 2130.35 ;
	END
END do27

PIN do26
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 1431.25 2129.1 1433.15 2130.35 ;
	END
END do26

PIN do25
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 1385.55 2129.1 1387.45 2130.35 ;
	END
END do25

PIN do24
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 1344.35 2129.1 1346.25 2130.35 ;
	END
END do24

PIN do23
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 1298.65 2129.1 1300.55 2130.35 ;
	END
END do23

PIN do22
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 1257.45 2129.1 1259.35 2130.35 ;
	END
END do22

PIN do21
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 1211.75 2129.1 1213.65 2130.35 ;
	END
END do21

PIN do20
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 1170.55 2129.1 1172.45 2130.35 ;
	END
END do20

PIN do19
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 1124.85 2129.1 1126.75 2130.35 ;
	END
END do19

PIN do18
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 1083.65 2129.1 1085.55 2130.35 ;
	END
END do18

PIN do17
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 1037.95 2129.1 1039.85 2130.35 ;
	END
END do17

PIN do16
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 996.75 2129.1 998.65 2130.35 ;
	END
END do16

PIN do15
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 951.05 2129.1 952.95 2130.35 ;
	END
END do15

PIN do14
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 909.85 2129.1 911.75 2130.35 ;
	END
END do14

PIN do13
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 864.15 2129.1 866.05 2130.35 ;
	END
END do13

PIN do12
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 822.95 2129.1 824.85 2130.35 ;
	END
END do12

PIN do11
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 777.25 2129.1 779.15 2130.35 ;
	END
END do11

PIN do10
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 736.05 2129.1 737.95 2130.35 ;
	END
END do10

PIN do9
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 690.35 2129.1 692.25 2130.35 ;
	END
END do9

PIN do8
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 649.16 2129.1 651.05 2130.35 ;
	END
END do8

PIN do7
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 603.45 2129.1 605.35 2130.35 ;
	END
END do7

PIN do6
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 562.25 2129.1 564.15 2130.35 ;
	END
END do6

PIN do5
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 516.55 2129.1 518.45 2130.35 ;
	END
END do5

PIN do4
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 475.35 2129.1 477.25 2130.35 ;
	END
END do4

PIN do3
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 429.65 2129.1 431.55 2130.35 ;
	END
END do3

PIN do2
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 388.45 2129.1 390.35 2130.35 ;
	END
END do2

PIN do1
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 342.75 2129.1 344.65 2130.35 ;
	END
END do1

PIN do0
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 301.55 2129.1 303.45 2130.35 ;
	END
END do0

PIN iwen3
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 1126.25 0.0 1128.25 1.25 ;
	END
END iwen3

PIN iwen2
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 1119.75 0.0 1121.75 1.25 ;
	END
END iwen2

PIN iwen1
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 1088.55 0.0 1090.55 1.25 ;
	END
END iwen1

PIN iwen0
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 1080.75 0.0 1082.75 1.25 ;
	END
END iwen0

PIN di31
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 1039.15 0.0 1041.15 1.25 ;
	END
END di31

PIN di30
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 1032.65 0.0 1034.65 1.25 ;
	END
END di30

PIN di29
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 1001.45 0.0 1003.45 1.25 ;
	END
END di29

PIN di28
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 993.65 0.0 995.65 1.25 ;
	END
END di28

PIN di27
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 952.05 0.0 954.05 1.25 ;
	END
END di27

PIN di26
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 945.55 0.0 947.55 1.25 ;
	END
END di26

PIN di25
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 914.35 0.0 916.35 1.25 ;
	END
END di25

PIN di24
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 907.85 0.0 909.85 1.25 ;
	END
END di24

PIN di23
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 866.25 0.0 868.25 1.25 ;
	END
END di23

PIN di22
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 858.45 0.0 860.45 1.25 ;
	END
END di22

PIN di21
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 827.25 0.0 829.25 1.25 ;
	END
END di21

PIN di20
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 820.75 0.0 822.75 1.25 ;
	END
END di20

PIN di19
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 779.15 0.0 781.15 1.25 ;
	END
END di19

PIN di18
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 771.35 0.0 773.35 1.25 ;
	END
END di18

PIN di17
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 740.15 0.0 742.15 1.25 ;
	END
END di17

PIN di16
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 733.65 0.0 735.65 1.25 ;
	END
END di16

PIN di15
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 692.05 0.0 694.05 1.25 ;
	END
END di15

PIN di14
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 684.25 0.0 686.25 1.25 ;
	END
END di14

PIN di13
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 654.35 0.0 656.35 1.25 ;
	END
END di13

PIN di12
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 646.55 0.0 648.55 1.25 ;
	END
END di12

PIN di11
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 604.95 0.0 606.95 1.25 ;
	END
END di11

PIN di10
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 597.15 0.0 599.15 1.25 ;
	END
END di10

PIN di9
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 567.25 0.0 569.25 1.25 ;
	END
END di9

PIN di8
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 559.45 0.0 561.45 1.25 ;
	END
END di8

PIN di7
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 517.85 0.0 519.85 1.25 ;
	END
END di7

PIN di6
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 511.35 0.0 513.35 1.25 ;
	END
END di6

PIN di5
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 480.15 0.0 482.15 1.25 ;
	END
END di5

PIN di4
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 472.35 0.0 474.35 1.25 ;
	END
END di4

PIN di3
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 430.75 0.0 432.75 1.25 ;
	END
END di3

PIN di2
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 424.25 0.0 426.25 1.25 ;
	END
END di2

PIN di1
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 393.05 0.0 395.05 1.25 ;
	END
END di1

PIN di0
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 385.25 0.0 387.25 1.25 ;
	END
END di0

PIN a0
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 161.65 0.0 163.65 1.25 ;
	END
END a0

PIN a1
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 144.75 0.0 146.75 1.25 ;
	END
END a1

PIN a2
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 134.35 0.0 136.35 1.25 ;
	END
END a2


PIN a3
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 93.75 0.0 95.75 1.25 ;
	END
END a3

PIN wrb
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 80.45 0.0 82.45 1.25 ;
	END
END wrb

PIN ceb
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 77.75 0.0 79.75 1.25 ;
	END
END ceb

PIN clk
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 66.75 0.0 68.75 1.25 ;
	END
END clk

PIN a4
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 59.35 0.0 61.35 1.25 ;
	END
END a4

PIN a5
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 55.95 0.0 57.95 1.25 ;
	END
END a5

PIN a6
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 51.15 0.0 53.15 1.25 ;
	END
END a6

PIN a7
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 42.05 0.0 44.05 1.25 ;
	END
END a7

PIN a8
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 36.85 0.0 38.85 1.25 ;
	END
END a8

PIN a9
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 27.75 0.0 29.75 1.25 ;
	END
END a9

PIN a10
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 22.55 0.0 24.55 1.25 ;
	END
END a10

	OBS
	LAYER Metal1 ;
RECT 1.40 1.40 1681.00 2128.95 ;
	LAYER Metal2 ;
RECT 1.40 1.40 1681.00 2128.95 ;
	LAYER Metal3 ;
RECT 1.40 1.40 1681.00 2128.95 ;
	LAYER Metal4 ;
RECT 1.40 1.40 1681.00 2128.95 ;
	END

END sram8k_pin
#1.12.03 u.j. + j.k. from GDS to lef

MACRO sram16k_pin
    CLASS BLOCK ;
    FOREIGN sram16k_pin 0 0 N ;
    SYMMETRY X Y r90 ;
    SIZE   1682.558 BY 3704.75 ;
    SITE core ;
    PIN vdd!
        USE power ;  
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT 1676.4 34.4 1682.4 65.65 ;
        RECT 1676.4 75.5 1682.4 81.75 ;
        RECT 1676.4 955.0 1682.4 961.25 ;
        RECT 1676.4 1845.0 1682.4 1851.25 ;
        RECT 1676.4 2736.25 1682.4 2742.5 ;
        RECT 1676.4 3622.15 1682.4 3628.4 ;
        RECT 1676.4 3638.75 1682.4 3670.0 ;
       RECT 0.0 3638.75 6.0 3670.0 ;
       RECT 0.0 3622.15 6.0 3628.4 ;
       RECT 0.0 2913.75 6.0 2920.0 ;
       RECT 0.0 2200.0 6.0 2206.25 ;
       RECT 0.0 1488.75 6.0 1495.0 ;
       RECT 0.0 775.0 6.0 781.25 ;
       RECT 0.0 75.5 6.0 81.75 ;
       RECT 0.0 34.4 6.0 65.65 ;
       END
    END vdd! 
    PIN vss!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ; 
        RECT 0.0 3671.25 6.0 3702.5 ;
        RECT 0.0 3629.65 6.0 3635.9 ;
        RECT 0.0 2921.25 6.0 2927.5 ;
        RECT 0.0 2207.5 6.0 2213.75 ;
        RECT 0.0 1496.25 6.0 1502.5 ;
        RECT 0.0 782.5 6.0 788.75 ;
        RECT 0.0 68.0 6.0 74.25 ;
        RECT 0.0 1.55 6.0 32.8 ;
        RECT 1676.4 1.55 1682.4 32.8 ;
        RECT 1676.4 68.0 1682.4 74.25 ;
        RECT 1676.4 962.5 1682.4 968.75 ;
        RECT 1676.4 1852.5 1682.4 1858.75 ;
        RECT 1676.4 2743.75 1682.4 2750.0 ;
        RECT 1676.4 3629.65 1682.4 3635.9 ;
        RECT 1676.4 3671.25 1682.4 3702.5 ;
        END
     END vss!



PIN oen3
	DIRECTION INPUT ;
	PORT
	LAYER Metal3 ;
	RECT 1328.15 3703.5 1330.15 3704.75 ;
	END
END oen3

PIN oen2
	DIRECTION INPUT ;
	PORT
	LAYER Metal3 ;
	RECT 980.55 3703.5 982.55 3704.75 ;
	END
END oen2

PIN oen1
	DIRECTION INPUT ;
	PORT
	LAYER Metal3 ;
	RECT 632.95 3703.5 634.95 3704.75 ;
	END
END oen1

PIN oen0
	DIRECTION INPUT ;
	PORT
	LAYER Metal3 ;
	RECT 285.35 3703.5 287.35 3704.75 ;
	END
END oen0

PIN do31
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 1646.2 3703.5 1648.2 3704.75 ;
	END
END do31

PIN do30
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 1605.0 3703.5 1607.0 3704.75 ;
	END
END do30

PIN do29
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 1559.3 3703.5 1561.3 3704.75 ;
	END
END do29

PIN do28
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 1518.1 3703.5 1520.1 3704.75 ;
	END
END do28

PIN do27
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 1472.4 3703.5 1474.4 3704.75 ;
	END
END do27

PIN do26
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 1431.2 3703.5 1433.2 3704.75 ;
	END
END do26

PIN do25
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 1385.5 3703.5 1387.5 3704.75 ;
	END
END do25

PIN do24
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 1344.3 3703.5 1346.3 3704.75 ;
	END
END do24

PIN do23
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 1298.6 3703.5 1300.6 3704.75 ;
	END
END do23

PIN do22
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 1257.4 3703.5 1259.4 3704.75 ;
	END
END do22

PIN do21
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 1211.7 3703.5 1213.7 3704.75 ;
	END
END do21

PIN do20
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 1170.5 3703.5 1172.5 3704.75 ;
	END
END do20

PIN do19
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 1124.8 3703.5 1126.8 3704.75 ;
	END
END do19

PIN do18
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 1083.6 3703.5 1085.6 3704.75 ;
	END
END do18

PIN do17
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 1037.9 3703.5 1039.9 3704.75 ;
	END
END do17

PIN do16
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 996.7 3703.5 998.7 3704.75 ;
	END
END do16

PIN do15
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 951.0 3703.5 953.0 3704.75 ;
	END
END do15

PIN do14
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 909.8 3703.5 911.8 3704.75 ;
	END
END do14

PIN do13
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 864.1 3703.5 866.1 3704.75 ;
	END
END do13

PIN do12
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 822.9 3703.5 824.9 3704.75 ;
	END
END do12

PIN do11
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 777.2 3703.5 779.2 3704.75 ;
	END
END do11

PIN do10
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 736.0 3703.5 738.0 3704.75 ;
	END
END do10

PIN do9
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 690.3 3703.5 692.3 3704.75 ;
	END
END do9

PIN do8
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 649.1 3703.5 651.1 3704.75 ;
	END
END do8

PIN do7
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 603.4 3703.5 605.4 3704.75 ;
	END
END do7

PIN do6
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 562.2 3703.5 564.2 3704.75 ;
	END
END do6

PIN do5
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 516.5 3703.5 518.5 3704.75 ;
	END
END do5

PIN do4
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 475.3 3703.5 477.3 3704.75 ;
	END
END do4

PIN do3
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 429.6 3703.5 431.6 3704.75 ;
	END
END do3

PIN do2
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 388.4 3703.5 390.4 3704.75 ;
	END
END do2

PIN do1
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 342.7 3703.5 344.7 3704.75 ;
	END
END do1

PIN do0
	DIRECTION OUTPUT ;
	PORT
	LAYER Metal2 ;
	RECT 301.5 3703.5 303.5 3704.75 ;
	END
END do0

PIN iwen3
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 1126.25 0.0 1128.25 1.25 ;
	END
END iwen3

PIN iwen2
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 1119.75 0.0 1121.75 1.25 ;
	END
END iwen2

PIN iwen1
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 1088.55 0.0 1090.55 1.25 ;
	END
END iwen1

PIN iwen0
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 1080.75 0.0 1082.75 1.25 ;
	END
END iwen0

PIN di31
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 1039.15 0.0 1041.15 1.25 ;
	END
END di31

PIN di30
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 1032.65 0.0 1034.65 1.25 ;
	END
END di30

PIN di29
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 1001.45 0.0 1003.45 1.25 ;
	END
END di29

PIN di28
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 993.65 0.0 995.65 1.25 ;
	END
END di28

PIN di27
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 952.05 0.0 954.05 1.25 ;
	END
END di27

PIN di26
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 945.55 0.0 947.55 1.25 ;
	END
END di26

PIN di25
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 914.35 0.0 916.35 1.25 ;
	END
END di25

PIN di24
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 907.85 0.0 909.85 1.25 ;
	END
END di24

PIN di23
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 866.25 0.0 868.25 1.25 ;
	END
END di23

PIN di22
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 858.45 0.0 860.45 1.25 ;
	END
END di22

PIN di21
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 827.25 0.0 829.25 1.25 ;
	END
END di21

PIN di20
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 820.75 0.0 822.75 1.25 ;
	END
END di20

PIN di19
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 779.15 0.0 781.15 1.25 ;
	END
END di19

PIN di18
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 771.35 0.0 773.35 1.25 ;
	END
END di18

PIN di17
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 740.15 0.0 742.15 1.25 ;
	END
END di17

PIN di16
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 733.65 0.0 735.65 1.25 ;
	END
END di16

PIN di15
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 692.05 0.0 694.05 1.25 ;
	END
END di15

PIN di14
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 684.25 0.0 686.25 1.25 ;
	END
END di14

PIN di13
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 654.35 0.0 656.35 1.25 ;
	END
END di13

PIN di12
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 646.55 0.0 648.55 1.25 ;
	END
END di12

PIN di11
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 604.95 0.0 606.95 1.25 ;
	END
END di11

PIN di10
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 597.15 0.0 599.15 1.25 ;
	END
END di10

PIN di9
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 567.25 0.0 569.25 1.25 ;
	END
END di9

PIN di8
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 559.45 0.0 561.45 1.25 ;
	END
END di8

PIN di7
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 517.85 0.0 519.85 1.25 ;
	END
END di7

PIN di6
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 511.35 0.0 513.35 1.25 ;
	END
END di6

PIN di5
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 480.15 0.0 482.15 1.25 ;
	END
END di5

PIN di4
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 472.35 0.0 474.35 1.25 ;
	END
END di4

PIN di3
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 430.75 0.0 432.75 1.25 ;
	END
END di3

PIN di2
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 424.25 0.0 426.25 1.25 ;
	END
END di2

PIN di1
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 393.05 0.0 395.05 1.25 ;
	END
END di1

PIN di0
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 385.25 0.0 387.25 1.25 ;
	END
END di0

PIN a0
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 161.65 0.0 163.65 1.25 ;
	END
END a0

PIN a1
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 144.75 0.0 146.75 1.25 ;
	END
END a1

PIN a2
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 134.35 0.0 136.35 1.25 ;
	END
END a2


PIN a3
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 93.75 0.0 95.75 1.25 ;
	END
END a3

PIN wrb
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 80.45 0.0 82.45 1.25 ;
	END
END wrb

PIN ceb
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 77.75 0.0 79.75 1.25 ;
	END
END ceb

PIN clk
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 66.75 0.0 68.75 1.25 ;
	END
END clk

PIN a4
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 59.35 0.0 61.35 1.25 ;
	END
END a4

PIN a5
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 55.95 0.0 57.95 1.25 ;
	END
END a5

PIN a6
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 51.15 0.0 53.15 1.25 ;
	END
END a6

PIN a7
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 42.05 0.0 44.05 1.25 ;
	END
END a7

PIN a8
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 36.85 0.0 38.85 1.25 ;
	END
END a8

PIN a9
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 27.75 0.0 29.75 1.25 ;
	END
END a9

PIN a10
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 22.55 0.0 24.55 1.25 ;
	END
END a10

PIN a11
	DIRECTION INPUT ;
	PORT
	LAYER Metal2 ;
	RECT 13.45 0.0 15.45 1.25 ;
	END
END a11
	OBS
	LAYER Metal1 ;
RECT 1.40 1.40 1681.00 3703.35 ;
	LAYER Metal2 ;
RECT 1.40 1.40 1681.00 3703.35 ;
	LAYER Metal3 ;
RECT 1.40 1.40 1681.00 3703.35 ;
	LAYER Metal4 ;
RECT 1.40 1.40 1681.00 3703.35 ;
	END

END sram16k_pin

#22.4.03 u.j. + j.k. from GDS to lef
#20.5.03 u.j. changed

#VERSION 5.4 ;

MACRO AFE
	CLASS BLOCK ;
	FOREIGN AFE 0 0 N ;
	SYMMETRY X Y ;
	SIZE  5510.00 BY 4723.75 ;
	SITE core ;

    PIN AGC_SEL 
        DIRECTION INPUT ; 
	PORT
	LAYER Metal4 ;
	RECT 5507.5 1202.5 5510.0 1205.0 ;
	END
    END AGC_SEL

    PIN RSSI 
        DIRECTION INPUT ; 
	PORT
	LAYER Metal4 ;
	RECT 5507.5 1197.5 5510.0 1200.0 ;
	END
    END RSSI

    PIN IF_AGC 
        DIRECTION INPUT ; 
	PORT
	LAYER Metal4 ;
	RECT 5507.5 1192.5 5510.0 1195.0 ;
	END
    END IF_AGC

    PIN LNA_GAIN 
        DIRECTION INPUT ; 
	PORT
	LAYER Metal4 ;
	RECT 5507.5 3917.45 5510.0 3919.95 ;
	END
    END LNA_GAIN

    PIN TX_GCi 
        DIRECTION INPUT ; 
	PORT
	LAYER Metal4 ;
	RECT 567.35 21.1 577.35 31.1 ;
	END
    END TX_GCi

    PIN TR_SW 
        DIRECTION INPUT ; 
	PORT
	LAYER Metal4 ;
	RECT 5507.5 3900.25 5510.0 3902.75 ;
	END
    END TR_SW

    PIN TX_Q 
        DIRECTION INPUT ; 
	PORT
	LAYER Metal4 ;
	RECT 1941.8 21.1 1951.8 31.1 ;
	END
    END TX_Q

    PIN TX_I 
        DIRECTION INPUT ; 
	PORT
	LAYER Metal4 ;
	RECT 1500.65 21.1 1510.65 31.1 ;
	END
    END TX_I

    PIN RX_In 
        DIRECTION OUTPUT ; 
	PORT
	LAYER Metal4 ;
	RECT 2794.05 21.1 2804.05 31.1 ;
	END
    END RX_In

    PIN RX_Ip 
        DIRECTION OUTPUT ; 
	PORT
	LAYER Metal4 ;
	RECT 2781.05 21.1 2791.05 31.1 ;
	END
    END RX_Ip

    PIN RX_Qn 
        DIRECTION OUTPUT ; 
	PORT
	LAYER Metal4 ;
	RECT 2341.9 21.1 2351.9 31.1 ;
	END
    END RX_Qn

    PIN RX_Qp 
        DIRECTION OUTPUT ; 
	PORT
	LAYER Metal4 ;
	RECT 2328.9 21.1 2338.9 31.1 ;
	END
    END RX_Qp

    PIN SYSCLK 
        DIRECTION INPUT ; 
	PORT
	LAYER Metal4 ;
	RECT 5507.5 3637.4 5510.0 3639.9 ;
	END
    END SYSCLK

    PIN RESET 
        DIRECTION INPUT ; 
	PORT
	LAYER Metal4 ;
	RECT 5507.5 3632.4 5510.0 3634.9 ;
	END
    END RESET

    PIN PLL_Set[0] 
        DIRECTION INPUT ; 
	PORT
	LAYER Metal4 ;
	RECT 5507.5 3627.4 5510.0 3629.9 ;
	END
    END PLL_Set[0]

    PIN PLL_Set[1] 
        DIRECTION INPUT ; 
	PORT
	LAYER Metal4 ;
	RECT 5507.5 3622.4 5510.0 3624.9 ;
	END
    END PLL_Set[1]

    PIN PLL_Set[2] 
        DIRECTION INPUT ; 
	PORT
	LAYER Metal4 ;
	RECT 5507.5 3617.4 5510.0 3619.9 ;
	END
    END PLL_Set[2]

    PIN PLL_Set[3] 
        DIRECTION INPUT ; 
	PORT
	LAYER Metal4 ;
	RECT 5507.5 3612.4 5510.0 3614.9 ;
	END
    END PLL_Set[3]

    PIN PLL_Set[4] 
        DIRECTION INPUT ; 
	PORT
	LAYER Metal4 ;
	RECT 5507.5 3607.4 5510.0 3609.9 ;
	END
    END PLL_Set[4]

    PIN PLL_Set[5] 
        DIRECTION INPUT ; 
	PORT
	LAYER Metal4 ;
	RECT 5507.5 3602.4 5510.0 3604.9 ;
	END
    END PLL_Set[5]

    PIN PLL_Set[6] 
        DIRECTION INPUT ; 
	PORT
	LAYER Metal4 ;
	RECT 5507.5 3597.4 5510.0 3599.9 ;
	END
    END PLL_Set[6]

    PIN PLL_Set[7] 
        DIRECTION INPUT ; 
	PORT
	LAYER Metal4 ;
	RECT 5507.5 3592.4 5510.0 3594.9 ;
	END
    END PLL_Set[7]

    PIN PLL_Set[8] 
        DIRECTION INPUT ; 
	PORT
	LAYER Metal4 ;
	RECT 5507.5 3587.4 5510.0 3589.9 ;
	END
    END PLL_Set[8]

    PIN PLL_Set[9] 
        DIRECTION INPUT ; 
	PORT
	LAYER Metal4 ;
	RECT 5507.5 3582.4 5510.0 3584.9 ;
	END
    END PLL_Set[9]

    PIN PLL_Set[10]
        DIRECTION INPUT ; 
	PORT
	LAYER Metal4 ;
	RECT 5507.5 3577.4 5510.0 3579.9 ;
	END
    END PLL_Set[10]

    PIN PLL_Set[11]
        DIRECTION INPUT ; 
	PORT
	LAYER Metal4 ;
	RECT 5507.5 3572.4 5510.0 3574.9 ;
	END
    END PLL_Set[11]

    PIN PLL_Set[12]
        DIRECTION INPUT ; 
	PORT
	LAYER Metal4 ;
	RECT 5507.5 3567.4 5510.0 3569.9 ;
	END
    END PLL_Set[12]

    PIN PLL_Set[13]
        DIRECTION INPUT ; 
	PORT
	LAYER Metal4 ;
	RECT 5507.5 3562.4 5510.0 3564.9 ;
	END
    END PLL_Set[13]

    PIN PLL_Set[14]
        DIRECTION INPUT ; 
	PORT
	LAYER Metal4 ;
	RECT 5507.5 3557.4 5510.0 3559.9 ;
	END
    END PLL_Set[14]

    PIN PLL_Set[15]
        DIRECTION INPUT ; 
	PORT
	LAYER Metal4 ;
	RECT 5507.5 3552.4 5510.0 3554.9 ;
	END
    END PLL_Set[15]

    PIN PLL_Set[16]
        DIRECTION INPUT ; 
	PORT
	LAYER Metal4 ;
	RECT 5507.5 3547.4 5510.0 3549.9 ;
	END
    END PLL_Set[16]

    PIN PLL_Set[17]
        DIRECTION INPUT ; 
	PORT
	LAYER Metal4 ;
	RECT 5507.5 3542.4 5510.0 3544.9 ;
	END
    END PLL_Set[17]

    PIN PLL_Set[18]
        DIRECTION INPUT ; 
	PORT
	LAYER Metal4 ;
	RECT 5507.5 3537.4 5510.0 3539.9 ;
	END
    END PLL_Set[18]

    PIN PLL_Set[19]
        DIRECTION INPUT ; 
	PORT
	LAYER Metal4 ;
	RECT 5507.5 3532.4 5510.0 3534.9 ;
	END
    END PLL_Set[19]
      OBS
        LAYER Metal1 ;
	RECT 0.00 31.10 5507.50 4723.75 ;
        LAYER Metal2 ;
	RECT 0.00 31.10 5507.50 4723.75 ;
        LAYER Metal3 ;
	RECT 0.00 31.10 5507.50 4723.75 ;
        LAYER Metal4 ;
	RECT 0.00 31.10 5507.50 4723.75 ;
        LAYER Metal5 ;
	RECT 0.00 31.10 5507.50 4723.75 ;
      END


END AFE
#24.04.03 + 11.06.03 u.j.

#VERSION 5.4 ;

MACRO RX_ADC
	CLASS BLOCK ;
	FOREIGN RX_ADC 0 0 N ;
	SYMMETRY X Y ;
	SIZE  1225.0 BY 1017.35 ;
	SITE core ;
    PIN vdd!
        USE power ;  
	DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal4 ;
        RECT  346.15 1013.05 352.95 1017.35 ;
        END
    END vdd!	
    PIN vss!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal4 ;	
        RECT 249.15 1012.25 257.0 1017.35 ;
        END
    END vss!	
    PIN vinvoltagen 
        DIRECTION INPUT ; 
	PORT
	LAYER Metal4 ;
	RECT 0.0 44.3 7.0 64.55 ;
	END
    END vinvoltagen
    PIN vinvoltagep 
        DIRECTION INPUT ; 
	PORT
	LAYER Metal4 ;
	RECT 0.0 237.4 4.2 242.5 ;
	END
    END vinvoltagep
    PIN mas_clk 
        DIRECTION INPUT ; 
	PORT
	LAYER Metal4 ;
	RECT 951.75 1015.6 954.25 1017.35 ;
	END
    END mas_clk
    PIN b[0] 
        DIRECTION OUTPUT ; 
	PORT
	LAYER Metal4 ;
	RECT 313.0 1014.95 315.5 1017.35 ;
	END
    END b[0]
    PIN b[1] 
        DIRECTION OUTPUT ; 
	PORT
	LAYER Metal4 ;
	RECT 393.0 1014.9 395.5 1017.35 ;
	END
    END b[1]
    PIN b[2] 
        DIRECTION OUTPUT ; 
	PORT
	LAYER Metal4 ;
	RECT 473.0 1014.95 475.5 1017.35 ;
	END
    END b[2]
    PIN b[3] 
        DIRECTION OUTPUT ; 
	PORT
	LAYER Metal4 ;
	RECT 553.0 1015.05 555.5 1017.35 ;
	END
    END b[3]
    PIN b[4] 
        DIRECTION OUTPUT ; 
	PORT
	LAYER Metal4 ;
	RECT 634.25 1015.2 636.75 1017.35 ;
	END
    END b[4]
    PIN b[5] 
        DIRECTION OUTPUT ; 
	PORT
	LAYER Metal4 ;
	RECT 713.0 1015.15 715.5 1017.35 ;
	END
    END b[5]
    PIN b[6] 
        DIRECTION OUTPUT ; 
	PORT
	LAYER Metal4 ;
	RECT 793.0 1015.15 795.5 1017.35 ;
	END
    END b[6]
    PIN b[7] 
        DIRECTION OUTPUT ; 
	PORT
	LAYER Metal4 ;
	RECT 874.25 1015.5 876.75 1017.35 ;
	END
    END b[7]
    PIN gnda! 
        USE ground ;
        DIRECTION INOUT ; 
	PORT
	LAYER Metal4 ;
	RECT 1216.6 5.05 1225.0 30.5 ;
	END
    END gnda!
    PIN vdda! 
        USE power ;  
        DIRECTION INOUT ; 
	PORT
	LAYER Metal4 ;
	RECT 1216.8 198.4 1224.8 279.2 ;
	END
    END vdda!
      OBS
        LAYER Metal1 ;
	RECT 4.0 2.0 1220.0 1015.6 ;
        LAYER Metal2 ;
	RECT 4.0 2.0 1220.0 1015.6 ;
        LAYER Metal3 ;
	RECT 4.0 2.0 1220.0 1015.6 ;
        LAYER Metal4 ;
	RECT 4.0 2.0 1220.0 1015.6 ;
      END
END RX_ADC

#24.04.03 11.06.03 u.j.

#VERSION 5.4 ;

MACRO RX_ADCSingle
	CLASS BLOCK ;
	FOREIGN RX_ADCSingle 0 0 N ;
	SYMMETRY X Y ;
	SIZE  1225.0 BY 1017.35 ;
	SITE core ;
    PIN vdd!
        USE power ;  
	DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal4 ;
        RECT  346.15 1013.05 352.95 1017.35 ;
        END
    END vdd!	
    PIN vss!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal4 ;	
        RECT 249.15 1012.25 257.0 1017.35 ;
        END
    END vss!	
    PIN vin 
        DIRECTION INPUT ; 
	PORT
	LAYER Metal4 ;
	RECT 0.0 44.3 7.0 64.55 ;
	END
    END vin
    PIN mas_clk 
        DIRECTION INPUT ; 
	PORT
	LAYER Metal4 ;
	RECT 951.75 1015.6 954.25 1017.35 ;
	END
    END mas_clk
    PIN b[0] 
        DIRECTION OUTPUT ; 
	PORT
	LAYER Metal4 ;
	RECT 313.0 1014.95 315.5 1017.35 ;
	END
    END b[0]
    PIN b[1] 
        DIRECTION OUTPUT ; 
	PORT
	LAYER Metal4 ;
	RECT 393.0 1014.9 395.5 1017.35 ;
	END
    END b[1]
    PIN b[2] 
        DIRECTION OUTPUT ; 
	PORT
	LAYER Metal4 ;
	RECT 473.0 1014.95 475.5 1017.35 ;
	END
    END b[2]
    PIN b[3] 
        DIRECTION OUTPUT ; 
	PORT
	LAYER Metal4 ;
	RECT 553.0 1015.05 555.5 1017.35 ;
	END
    END b[3]
    PIN b[4] 
        DIRECTION OUTPUT ; 
	PORT
	LAYER Metal4 ;
	RECT 634.25 1015.2 636.75 1017.35 ;
	END
    END b[4]
    PIN b[5] 
        DIRECTION OUTPUT ; 
	PORT
	LAYER Metal4 ;
	RECT 713.0 1015.15 715.5 1017.35 ;
	END
    END b[5]
    PIN b[6] 
        DIRECTION OUTPUT ; 
	PORT
	LAYER Metal4 ;
	RECT 793.0 1015.15 795.5 1017.35 ;
	END
    END b[6]
    PIN b[7] 
        DIRECTION OUTPUT ; 
	PORT
	LAYER Metal4 ;
	RECT 874.25 1015.5 876.75 1017.35 ;
	END
    END b[7]
    PIN gnda! 
        USE ground ;
        DIRECTION INOUT ; 
	PORT
	LAYER Metal4 ;
	RECT 1216.6 5.05 1225.0 30.5 ;
	END
    END gnda!
    PIN vdda! 
        USE power ;  
        DIRECTION INOUT ; 
	PORT
	LAYER Metal4 ;
	RECT 1216.8 198.4 1224.8 279.2 ;
	END
    END vdda!
      OBS
        LAYER Metal1 ;
	RECT 4.0 2.0 1220.0 1015.6 ;
        LAYER Metal2 ;
	RECT 4.0 2.0 1220.0 1015.6 ;
        LAYER Metal3 ;
	RECT 4.0 2.0 1220.0 1015.6 ;
        LAYER Metal4 ;
	RECT 4.0 2.0 1220.0 1015.6 ;
      END
END RX_ADCSingle


#24.04.03 u.j. 22.05.03

#VERSION 5.4 ;

MACRO TX_DAC
	CLASS BLOCK ;
	FOREIGN TX_DAC 0 0 N ;
	SYMMETRY X Y ;
	SIZE  1108.0 BY 1050.0 ;
	SITE core ;
    PIN vdd!
        USE power ;  
	DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal4 ;
        RECT  162.65 1045.1 172.65 1050.0 ;
        END
    END vdd!	
    PIN vss!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal4 ;	
        RECT 882.5 1042.9 912.5 1049.8 ;
        END
    END vss!	

    PIN Clock 
        DIRECTION INPUT ; 
	PORT
	LAYER Metal4 ;
	RECT 743.4 1048.1 745.9 1050.0 ;
	END
    END Clock
    PIN TX_DATA[0] 
        DIRECTION INPUT ; 
	PORT
	LAYER Metal4 ;
	RECT 213.95 1047.85 216.45 1050.0 ;
	END
    END TX_DATA[0]
    PIN TX_DATA[1] 
        DIRECTION INPUT ; 
	PORT
	LAYER Metal4 ;
	RECT 256.4 1048.6 258.9 1050.0 ;
	END
    END TX_DATA[1]
    PIN TX_DATA[2] 
        DIRECTION INPUT ; 
	PORT
	LAYER Metal4 ;
	RECT 308.9 1048.75 311.4 1050.0 ;
	END
    END TX_DATA[2]
    PIN TX_DATA[3] 
        DIRECTION INPUT ; 
	PORT
	LAYER Metal4 ;
	RECT 362.65 1048.35 365.15 1050.0 ;
	END
    END TX_DATA[3]
    PIN TX_DATA[4] 
        DIRECTION INPUT ; 
	PORT
	LAYER Metal4 ;
	RECT 415.85 1048.35 418.35 1050.0 ;
	END
    END TX_DATA[4]
    PIN TX_DATA[5] 
        DIRECTION INPUT ; 
	PORT
	LAYER Metal4 ;
	RECT 470.1 1048.35 472.6 1050.0 ;
	END
    END TX_DATA[5]
    PIN TX_DATA[6] 
        DIRECTION INPUT ; 
	PORT
	LAYER Metal4 ;
	RECT 525.2 1048.45 527.7 1049.95 ;
	END
    END TX_DATA[6]
    PIN TX_DATA[7] 
        DIRECTION INPUT ; 
	PORT
	LAYER Metal4 ;
	RECT 579.05 1048.3 581.55 1050.0 ;
	END
    END TX_DATA[7]
    PIN TX_DATA[8] 
        DIRECTION INPUT ; 
	PORT
	LAYER Metal4 ;
	RECT 635.2 1048.1 637.65 1050.0 ;
	END
    END TX_DATA[8]
    PIN TX_DATA[9] 
        DIRECTION INPUT ; 
	PORT
	LAYER Metal4 ;
	RECT 687.65 1048.75 691.4 1050.0 ;
	END
    END TX_DATA[9]
    PIN DAC_OP 
        DIRECTION OUTPUT ; 
	PORT
	LAYER Metal4 ;
	RECT 1095.5 99.1 1107.4 150.3 ;
	END
    END DAC_OP
    PIN gnda! 
        USE ground ;
        DIRECTION INOUT ; 
	PORT
	LAYER Metal4 ;
	RECT 1097.5 2.5 1107.4 57.9 ;
	END
    END gnda!
    PIN vdda! 
        USE power ;  
        DIRECTION INOUT ; 
	PORT
	LAYER Metal4 ;
	RECT 1094.8 252.2 1107.3 314.3 ;
	END
    END vdda!
      OBS
        LAYER Metal1 ;
	RECT 0.00 0.00 1103.00 1048.00 ;
        LAYER Metal2 ;
	RECT 0.00 0.00 1103.00 1048.00 ;
        LAYER Metal3 ;
	RECT 0.00 0.00 1103.00 1048.00 ;
        LAYER Metal4 ;
	RECT 0.00 0.00 1103.00 1048.00 ;
      END
END TX_DAC


#24.04.03 u.j. 22.05.03
VERSION 5.4 ;
MACRO TX_DACSingle
	CLASS BLOCK ;
	FOREIGN TX_DACSingle 0 0 N ;
	SYMMETRY X Y ;
	SIZE  600.0 BY 600.0 ;
	SITE core ;
    PIN vdd!
        USE power ;  
	DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal4 ;
        RECT  156.15 589.8 184.9 600.0 ;
        END
    END vdd!	
    PIN vss!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal4 ;	
        RECT 79.05 592.9 90.0 600.0 ;
        END
    END vss!	

    PIN Clock 
        DIRECTION INPUT ; 
	PORT
	LAYER Metal4 ;
	RECT 431.9 598.8 434.4 600.0 ;
	END
    END Clock
    PIN TX_DATA[0] 
        DIRECTION INPUT ; 
	PORT
	LAYER Metal4 ;
	RECT 234.4 598.5 236.9 600.0 ;
	END
    END TX_DATA[0]
    PIN TX_DATA[1] 
        DIRECTION INPUT ; 
	PORT
	LAYER Metal4 ;
	RECT 259.4 598.25 261.9 600.0 ;
	END
    END TX_DATA[1]
    PIN TX_DATA[2] 
        DIRECTION INPUT ; 
	PORT
	LAYER Metal4 ;
	RECT 283.15 598.15 285.65 600.0 ;
	END
    END TX_DATA[2]
    PIN TX_DATA[3] 
        DIRECTION INPUT ; 
	PORT
	LAYER Metal4 ;
	RECT 309.4 598.2 311.9 600.0 ;
	END
    END TX_DATA[3]
    PIN TX_DATA[4] 
        DIRECTION INPUT ; 
	PORT
	LAYER Metal4 ;
	RECT 334.4 598.75 336.9 600.0 ;
	END
    END TX_DATA[4]
    PIN TX_DATA[5] 
        DIRECTION INPUT ; 
	PORT
	LAYER Metal4 ;
	RECT 359.4 598.75 361.9 600.0 ;
	END
    END TX_DATA[5]
    PIN TX_DATA[6] 
        DIRECTION INPUT ; 
	PORT
	LAYER Metal4 ;
	RECT 384.4 598.15 386.9 600.0 ;
	END
    END TX_DATA[6]
    PIN TX_DATA[7] 
        DIRECTION INPUT ; 
	PORT
	LAYER Metal4 ;
	RECT 409.4 598.35 411.9 600.0 ;
	END
    END TX_DATA[7]
    PIN DAC_OP 
        DIRECTION OUTPUT ; 
	PORT
	LAYER Metal4 ;
	RECT 592.45 104.1 600.0 126.15 ;
	END
    END DAC_OP
    PIN gnda! 
        USE ground ;
        DIRECTION INOUT ; 
	PORT
	LAYER Metal4 ;
	RECT 591.5 32.9 600.0 52.45 ;
	END
    END gnda!
    PIN vdda! 
        USE power ;  
        DIRECTION INOUT ; 
	PORT
	LAYER Metal4 ;
	RECT 596.15 167.9 600.0 202.15 ;
	END
    END vdda!
      OBS
        LAYER Metal1 ;
	RECT 0.00 0.00 597.00 598.50 ;
        LAYER Metal2 ;
	RECT 0.00 0.00 597.00 598.50 ;
        LAYER Metal3 ;
	RECT 0.00 0.00 597.00 598.50 ;
        LAYER Metal4 ;
	RECT 0.00 0.00 597.00 598.50 ;
      END
END TX_DACSingle


MACRO GSRAMm128_128_32dbf
  CLASS BLOCK ;
  FOREIGN GSRAMm128_128_32dbf  0 0 N ;
  SIZE 987.00 BY 1354.80 ;
  SYMMETRY x y r90 ;
  SITE core ;
  PIN ADR[6]
    DIRECTION INPUT ;
    PORT 
    LAYER Metal1 ;
    RECT  74.60 1340.80 75.40 1341.80 ;
  END
  END ADR[6]
  PIN ADR[5]
    DIRECTION INPUT ;
    PORT 
    LAYER Metal1 ;
    RECT  86.500  1340.800  87.300  1341.800 ;
    END
  END ADR[5]
  PIN ADR[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.015 ;
    PORT 
      LAYER Metal1 ;
        RECT  98.400  1340.800  99.200  1341.800 ;
    END
  END ADR[4]
  PIN ADR[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.015 ;
    PORT 
      LAYER Metal1 ;
        RECT  110.300  1340.800  111.100  1341.800 ;
    END
  END ADR[3]
  PIN ADR[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.015 ;
    PORT 
      LAYER Metal1 ;
        RECT  122.200  1340.800  123.000  1341.800 ;
    END
  END ADR[2]
  PIN ADR[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.015 ;
    PORT 
      LAYER Metal1 ;
        RECT  134.100  1340.800  134.900  1341.800 ;
    END
  END ADR[1]
  PIN ADR[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.015 ;
    PORT 
      LAYER Metal1 ;
        RECT  146.000  1340.800  146.800  1341.800 ;
    END
  END ADR[0]
  PIN RDSTR
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.015 ;
    PORT 
      LAYER Metal3 ;
        RECT  -1.000  368.400  0.000  370.300 ;
    END
  END RDSTR
  PIN WRSTR
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.015 ;
    PORT 
      LAYER Metal3 ;
        RECT  -1.000  363.900  0.000  365.800 ;
    END
  END WRSTR
  PIN MASK[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.015 ;
    PORT 
      LAYER Metal3 ;
        RECT  -1.000  351.450  0.000  352.050 ;
    END
  END MASK[0]
  PIN MASK[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.015 ;
    PORT 
      LAYER Metal3 ;
        RECT  -1.000  352.700  0.000  353.300 ;
    END
  END MASK[1]
  PIN MASK[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.015 ;
    PORT 
      LAYER Metal3 ;
        RECT  -1.000  353.950  0.000  354.550 ;
    END
  END MASK[2]
  PIN MASK[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.015 ;
    PORT 
      LAYER Metal3 ;
        RECT  -1.000  355.200  0.000  355.800 ;
    END
  END MASK[3]
  PIN CS
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.015 ;
    PORT 
      LAYER Metal3 ;
        RECT  -1.000  357.200  0.000  359.100 ;
    END
  END CS
  PIN STOP
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.001 ;
    PORT 
      LAYER Metal1 ;
        RECT  215.550  -1.000  216.350  0.000 ;
    END
  END STOP
  PIN BIST
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.023 ;
    PORT 
      LAYER Metal1 ;
        RECT  254.850  -1.000  255.650  0.000 ;
    END
  END BIST
  PIN COMP_OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.001 ;
    PORT 
      LAYER Metal3 ;
        RECT  987.000  126.150  988.000  126.750 ;
    END
  END COMP_OUT
  PIN OUT[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.001 ;
    PORT 
      LAYER Metal1 ;
        RECT  261.000  -1.000  264.000  0.000 ;
    END
  END OUT[0]
  PIN OUT[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.001 ;
    PORT 
      LAYER Metal1 ;
        RECT  281.200  -1.000  284.200  0.000 ;
    END
  END OUT[1]
  PIN OUT[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.001 ;
    PORT 
      LAYER Metal1 ;
        RECT  301.400  -1.000  304.400  0.000 ;
    END
  END OUT[2]
  PIN OUT[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.001 ;
    PORT 
      LAYER Metal1 ;
        RECT  321.600  -1.000  324.600  0.000 ;
    END
  END OUT[3]
  PIN OUT[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.001 ;
    PORT 
      LAYER Metal1 ;
        RECT  345.450  -1.000  348.450  0.000 ;
    END
  END OUT[4]
  PIN OUT[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.001 ;
    PORT 
      LAYER Metal1 ;
        RECT  365.650  -1.000  368.650  0.000 ;
    END
  END OUT[5]
  PIN OUT[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.001 ;
    PORT 
      LAYER Metal1 ;
        RECT  385.850  -1.000  388.850  0.000 ;
    END
  END OUT[6]
  PIN OUT[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.001 ;
    PORT 
      LAYER Metal1 ;
        RECT  406.050  -1.000  409.050  0.000 ;
    END
  END OUT[7]
  PIN OUT[8]
    DIRECTION OUTPUT ;
    PORT 
      LAYER Metal1 ;
        RECT  429.900  -1.000  432.900  0.000 ;
    END
  END OUT[8]
  PIN OUT[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.001 ;
    PORT 
      LAYER Metal1 ;
        RECT  450.100  -1.000  453.100  0.000 ;
    END
  END OUT[9]
  PIN OUT[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.001 ;
    PORT 
      LAYER Metal1 ;
        RECT  470.300  -1.000  473.300  0.000 ;
    END
  END OUT[10]
  PIN OUT[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.001 ;
    PORT 
      LAYER Metal1 ;
        RECT  490.500  -1.000  493.500  0.000 ;
    END
  END OUT[11]
  PIN OUT[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.001 ;
    PORT 
      LAYER Metal1 ;
        RECT  514.350  -1.000  517.350  0.000 ;
    END
  END OUT[12]
  PIN OUT[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.001 ;
    PORT 
      LAYER Metal1 ;
        RECT  534.550  -1.000  537.550  0.000 ;
    END
  END OUT[13]
  PIN OUT[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.001 ;
    PORT 
      LAYER Metal1 ;
        RECT  554.750  -1.000  557.750  0.000 ;
    END
  END OUT[14]
  PIN OUT[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.001 ;
    PORT 
      LAYER Metal1 ;
        RECT  574.950  -1.000  577.950  0.000 ;
    END
  END OUT[15]
  PIN OUT[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.001 ;
    PORT 
      LAYER Metal1 ;
        RECT  598.800  -1.000  601.800  0.000 ;
    END
  END OUT[16]
  PIN OUT[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.001 ;
    PORT 
      LAYER Metal1 ;
        RECT  619.000  -1.000  622.000  0.000 ;
    END
  END OUT[17]
  PIN OUT[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.001 ;
    PORT 
      LAYER Metal1 ;
        RECT  639.200  -1.000  642.200  0.000 ;
    END
  END OUT[18]
  PIN OUT[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.001 ;
    PORT 
      LAYER Metal1 ;
        RECT  659.400  -1.000  662.400  0.000 ;
    END
  END OUT[19]
  PIN OUT[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.001 ;
    PORT 
      LAYER Metal1 ;
        RECT  683.250  -1.000  686.250  0.000 ;
    END
  END OUT[20]
  PIN OUT[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.001 ;
    PORT 
      LAYER Metal1 ;
        RECT  703.450  -1.000  706.450  0.000 ;
    END
  END OUT[21]
  PIN OUT[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.001 ;
    PORT 
      LAYER Metal1 ;
        RECT  723.650  -1.000  726.650  0.000 ;
    END
  END OUT[22]
  PIN OUT[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.001 ;
    PORT 
      LAYER Metal1 ;
        RECT  743.850  -1.000  746.850  0.000 ;
    END
  END OUT[23]
  PIN OUT[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.001 ;
    PORT 
      LAYER Metal1 ;
        RECT  767.700  -1.000  770.700  0.000 ;
    END
  END OUT[24]
  PIN OUT[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.001 ;
    PORT 
      LAYER Metal1 ;
        RECT  787.900  -1.000  790.900  0.000 ;
    END
  END OUT[25]
  PIN OUT[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.001 ;
    PORT 
      LAYER Metal1 ;
        RECT  808.100  -1.000  811.100  0.000 ;
    END
  END OUT[26]
  PIN OUT[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.001 ;
    PORT 
      LAYER Metal1 ;
        RECT  828.300  -1.000  831.300  0.000 ;
    END
  END OUT[27]
  PIN OUT[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.001 ;
    PORT 
      LAYER Metal1 ;
        RECT  852.150  -1.000  855.150  0.000 ;
    END
  END OUT[28]
  PIN OUT[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.001 ;
    PORT 
      LAYER Metal1 ;
        RECT  872.350  -1.000  875.350  0.000 ;
    END
  END OUT[29]
  PIN OUT[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.001 ;
    PORT 
      LAYER Metal1 ;
        RECT  892.550  -1.000  895.550  0.000 ;
    END
  END OUT[30]
  PIN OUT[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.001 ;
    PORT 
      LAYER Metal1 ;
        RECT  912.750  -1.000  915.750  0.000 ;
    END
  END OUT[31]
  PIN DATA[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.007 ;
    PORT 
      LAYER Metal1 ;
        RECT  252.500  -1.000  253.500  0.000 ;
    END
  END DATA[0]
  PIN DATA[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.007 ;
    PORT 
      LAYER Metal1 ;
        RECT  272.700  -1.000  273.700  0.000 ;
    END
  END DATA[1]
  PIN DATA[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.007 ;
    PORT 
      LAYER Metal1 ;
        RECT  292.900  -1.000  293.900  0.000 ;
    END
  END DATA[2]
  PIN DATA[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.007 ;
    PORT 
      LAYER Metal1 ;
        RECT  313.100  -1.000  314.100  0.000 ;
    END
  END DATA[3]
  PIN DATA[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.007 ;
    PORT 
      LAYER Metal1 ;
        RECT  336.950  -1.000  337.950  0.000 ;
    END
  END DATA[4]
  PIN DATA[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.007 ;
    PORT 
      LAYER Metal1 ;
        RECT  357.150  -1.000  358.150  0.000 ;
    END
  END DATA[5]
  PIN DATA[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.007 ;
    PORT 
      LAYER Metal1 ;
        RECT  377.350  -1.000  378.350  0.000 ;
    END
  END DATA[6]
  PIN DATA[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.007 ;
    PORT 
      LAYER Metal1 ;
        RECT  397.550  -1.000  398.550  0.000 ;
    END
  END DATA[7]
  PIN DATA[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.007 ;
    PORT 
      LAYER Metal1 ;
        RECT  421.400  -1.000  422.400  0.000 ;
    END
  END DATA[8]
  PIN DATA[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.007 ;
    PORT 
      LAYER Metal1 ;
        RECT  441.600  -1.000  442.600  0.000 ;
    END
  END DATA[9]
  PIN DATA[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.007 ;
    PORT 
      LAYER Metal1 ;
        RECT  461.800  -1.000  462.800  0.000 ;
    END
  END DATA[10]
  PIN DATA[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.007 ;
    PORT 
      LAYER Metal1 ;
        RECT  482.000  -1.000  483.000  0.000 ;
    END
  END DATA[11]
  PIN DATA[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.007 ;
    PORT 
      LAYER Metal1 ;
        RECT  505.850  -1.000  506.850  0.000 ;
    END
  END DATA[12]
  PIN DATA[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.007 ;
    PORT 
      LAYER Metal1 ;
        RECT  526.050  -1.000  527.050  0.000 ;
    END
  END DATA[13]
  PIN DATA[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.007 ;
    PORT 
      LAYER Metal1 ;
        RECT  546.250  -1.000  547.250  0.000 ;
    END
  END DATA[14]
  PIN DATA[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.007 ;
    PORT 
      LAYER Metal1 ;
        RECT  566.450  -1.000  567.450  0.000 ;
    END
  END DATA[15]
  PIN DATA[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.007 ;
    PORT 
      LAYER Metal1 ;
        RECT  590.300  -1.000  591.300  0.000 ;
    END
  END DATA[16]
  PIN DATA[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.007 ;
    PORT 
      LAYER Metal1 ;
        RECT  610.500  -1.000  611.500  0.000 ;
    END
  END DATA[17]
  PIN DATA[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.007 ;
    PORT 
      LAYER Metal1 ;
        RECT  630.700  -1.000  631.700  0.000 ;
    END
  END DATA[18]
  PIN DATA[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.007 ;
    PORT 
      LAYER Metal1 ;
        RECT  650.900  -1.000  651.900  0.000 ;
    END
  END DATA[19]
  PIN DATA[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.007 ;
    PORT 
      LAYER Metal1 ;
        RECT  674.750  -1.000  675.750  0.000 ;
    END
  END DATA[20]
  PIN DATA[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.007 ;
    PORT 
      LAYER Metal1 ;
        RECT  694.950  -1.000  695.950  0.000 ;
    END
  END DATA[21]
  PIN DATA[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.007 ;
    PORT 
      LAYER Metal1 ;
        RECT  715.150  -1.000  716.150  0.000 ;
    END
  END DATA[22]
  PIN DATA[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.007 ;
    PORT 
      LAYER Metal1 ;
        RECT  735.350  -1.000  736.350  0.000 ;
    END
  END DATA[23]
  PIN DATA[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.007 ;
    PORT 
      LAYER Metal1 ;
        RECT  759.200  -1.000  760.200  0.000 ;
    END
  END DATA[24]
  PIN DATA[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.007 ;
    PORT 
      LAYER Metal1 ;
        RECT  779.400  -1.000  780.400  0.000 ;
    END
  END DATA[25]
  PIN DATA[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.007 ;
    PORT 
      LAYER Metal1 ;
        RECT  799.600  -1.000  800.600  0.000 ;
    END
  END DATA[26]
  PIN DATA[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    CAPACITANCE 0.007 ;
    PORT 
      LAYER Metal1 ;
        RECT  819.800  -1.000  820.800  0.000 ;
    END
  END DATA[27]
  PIN DATA[28]
    DIRECTION INPUT ;
    PORT 
      LAYER Metal1 ;
        RECT  843.650  -1.000  844.650  0.000 ;
    END
  END DATA[28]
  PIN DATA[29]
    DIRECTION INPUT ;
    PORT 
      LAYER Metal1 ;
        RECT  863.850  -1.000  864.850  0.000 ;
    END
  END DATA[29]
  PIN DATA[30]
    DIRECTION INPUT ;
    PORT 
      LAYER Metal1 ;
        RECT  884.050  -1.000  885.050  0.000 ;
    END
  END DATA[30]
  PIN DATA[31]
    DIRECTION INPUT ;
    PORT 
      LAYER Metal1 ;
        RECT  904.250  -1.000  905.250  0.000 ;
    END
  END DATA[31]
  PIN ADR[7]
    DIRECTION INPUT ;
    PORT 
      LAYER Metal3 ;
        RECT  -1.000  240.600  0.000  241.200 ;
    END
  END ADR[7]
  PIN ADR[8]
    DIRECTION INPUT ;
    PORT 
      LAYER Metal3 ;
        RECT  -1.000  238.100  0.000  238.700 ;
    END
  END ADR[8]
  PIN CLK
    PORT    
      LAYER Metal3 ;
        RECT  -1.000  373.950  0.000  379.950 ;
    END
  END CLK
    PIN vdd!
        USE power ;  
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal1 ;
        RECT  32.000  1324.800  62.000  1354.800 ;
        RECT  925.000  1324.800  955.000  1354.800 ;
        RECT  32.000  0.000  62.000  30.000 ;
        RECT  925.000  0.000  955.000  30.000 ;
    END
  END vdd!
   PIN vss!
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER Metal2 ; 
        RECT  32.000  1324.800  62.000  1354.800 ;
        RECT  925.000  1324.800  955.000  1354.800 ;
        RECT  32.000  0.000  62.000  30.000 ;
        RECT  925.000  0.000  955.000  30.000 ;
    END
  END vss!
  OBS
    LAYER Metal1 ;
      RECT  51.000  0.000  955.000  1340.800 ;
    LAYER Metal2 ;
      RECT  0.000  0.000  987.000  1354.800 ;
    LAYER Metal3 ;
      RECT  0.000  67.000  987.000  1276.800 ;
  END
END GSRAMm128_128_32dbf
END LIBRARY
